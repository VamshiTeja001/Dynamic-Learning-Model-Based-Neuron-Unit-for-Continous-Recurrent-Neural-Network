
`timescale 1ns / 1ps


//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 25.02.2025 00:56:53
// Design Name: 
// Module Name: Sigmoid
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Sigmoid(
input [31:0] numb,
input rst,
input clk,
output reg [31:0] sigmoid_out


    );
    
    reg x =0;
    
    reg [7:0] exponent;
    reg [22:0] mantissa;
    reg sign;
    real float_value,scaled_value, rounded_value;
    reg [31:0] result;
    integer int_scaled_value;
    always @(*) begin
        // Extract sign, exponent, and mantissa
        sign = numb[31];
        exponent = numb[30:23];
        mantissa = numb[22:0];

        // Convert IEEE 754 to floating-point value
        float_value = (1.0 + (mantissa / (2**23))) * (2**(exponent - 127));
        if (sign == 1) float_value = -float_value;

      // Scale by 100
        scaled_value = float_value * 100.0;
        
        // Convert to integer (truncating the decimal)
        int_scaled_value = scaled_value;  // Implicit truncation of decimal part

        // Convert back to real (divide by 100)
        rounded_value = int_scaled_value / 100.0;

        // Convert back to IEEE 754
        sign = (rounded_value < 0) ? 1 : 0;
        if (sign) rounded_value = -rounded_value;

        exponent = 127;
        while (rounded_value >= 2.0) begin
            rounded_value = rounded_value / 2.0;
            exponent = exponent + 1;
        end
        while (rounded_value < 1.0 && rounded_value != 0.0) begin
            rounded_value = rounded_value * 2.0;
            exponent = exponent - 1;
        end

        mantissa = (rounded_value - 1.0) * (2**23);

        // Construct IEEE 754 output
        x = {sign, exponent, mantissa};
        end
    
    always@(posedge clk or posedge rst)
begin
if (rst) sigmoid_out=0;
else begin

//case(x)
case (numb)
        32'hC0C00000: sigmoid_out = 32'h3B220BBC; // -6.00 -> sigmoid(-6.00) = 0.00247262
        32'hC0BFAE14: sigmoid_out = 32'h3B23AB9C; // -5.99 -> sigmoid(-5.99) = 0.00249741
        32'hC0BF5C29: sigmoid_out = 32'h3B254FA5; // -5.98 -> sigmoid(-5.98) = 0.00252245
        32'hC0BF0A3D: sigmoid_out = 32'h3B26F7E2; // -5.97 -> sigmoid(-5.97) = 0.00254773
        32'hC0BEB852: sigmoid_out = 32'h3B28A45C; // -5.96 -> sigmoid(-5.96) = 0.00257327
        32'hC0BE6666: sigmoid_out = 32'h3B2A551F; // -5.95 -> sigmoid(-5.95) = 0.00259907
        32'hC0BE147B: sigmoid_out = 32'h3B2C0A36; // -5.94 -> sigmoid(-5.94) = 0.00262512
        32'hC0BDC28F: sigmoid_out = 32'h3B2DC3AB; // -5.93 -> sigmoid(-5.93) = 0.00265143
        32'hC0BD70A4: sigmoid_out = 32'h3B2F818A; // -5.92 -> sigmoid(-5.92) = 0.00267801
        32'hC0BD1EB8: sigmoid_out = 32'h3B3143DE; // -5.91 -> sigmoid(-5.91) = 0.00270485
        32'hC0BCCCCD: sigmoid_out = 32'h3B330AB2; // -5.90 -> sigmoid(-5.90) = 0.00273196
        32'hC0BC7AE1: sigmoid_out = 32'h3B34D612; // -5.89 -> sigmoid(-5.89) = 0.00275934
        32'hC0BC28F6: sigmoid_out = 32'h3B36A60A; // -5.88 -> sigmoid(-5.88) = 0.00278700
        32'hC0BBD70A: sigmoid_out = 32'h3B387AA4; // -5.87 -> sigmoid(-5.87) = 0.00281493
        32'hC0BB851F: sigmoid_out = 32'h3B3A53ED; // -5.86 -> sigmoid(-5.86) = 0.00284314
        32'hC0BB3333: sigmoid_out = 32'h3B3C31F1; // -5.85 -> sigmoid(-5.85) = 0.00287163
        32'hC0BAE148: sigmoid_out = 32'h3B3E14BC; // -5.84 -> sigmoid(-5.84) = 0.00290041
        32'hC0BA8F5C: sigmoid_out = 32'h3B3FFC5A; // -5.83 -> sigmoid(-5.83) = 0.00292947
        32'hC0BA3D71: sigmoid_out = 32'h3B41E8D7; // -5.82 -> sigmoid(-5.82) = 0.00295882
        32'hC0B9EB85: sigmoid_out = 32'h3B43DA3F; // -5.81 -> sigmoid(-5.81) = 0.00298847
        32'hC0B9999A: sigmoid_out = 32'h3B45D09F; // -5.80 -> sigmoid(-5.80) = 0.00301842
        32'hC0B947AE: sigmoid_out = 32'h3B47CC05; // -5.79 -> sigmoid(-5.79) = 0.00304866
        32'hC0B8F5C3: sigmoid_out = 32'h3B49CC7B; // -5.78 -> sigmoid(-5.78) = 0.00307920
        32'hC0B8A3D7: sigmoid_out = 32'h3B4BD210; // -5.77 -> sigmoid(-5.77) = 0.00311005
        32'hC0B851EC: sigmoid_out = 32'h3B4DDCD0; // -5.76 -> sigmoid(-5.76) = 0.00314121
        32'hC0B80000: sigmoid_out = 32'h3B4FECC9; // -5.75 -> sigmoid(-5.75) = 0.00317268
        32'hC0B7AE14: sigmoid_out = 32'h3B520207; // -5.74 -> sigmoid(-5.74) = 0.00320447
        32'hC0B75C29: sigmoid_out = 32'h3B541C99; // -5.73 -> sigmoid(-5.73) = 0.00323657
        32'hC0B70A3D: sigmoid_out = 32'h3B563C8B; // -5.72 -> sigmoid(-5.72) = 0.00326899
        32'hC0B6B852: sigmoid_out = 32'h3B5861EC; // -5.71 -> sigmoid(-5.71) = 0.00330173
        32'hC0B66666: sigmoid_out = 32'h3B5A8CC8; // -5.70 -> sigmoid(-5.70) = 0.00333481
        32'hC0B6147B: sigmoid_out = 32'h3B5CBD2F; // -5.69 -> sigmoid(-5.69) = 0.00336821
        32'hC0B5C28F: sigmoid_out = 32'h3B5EF32E; // -5.68 -> sigmoid(-5.68) = 0.00340195
        32'hC0B570A4: sigmoid_out = 32'h3B612ED2; // -5.67 -> sigmoid(-5.67) = 0.00343602
        32'hC0B51EB8: sigmoid_out = 32'h3B63702C; // -5.66 -> sigmoid(-5.66) = 0.00347043
        32'hC0B4CCCD: sigmoid_out = 32'h3B65B748; // -5.65 -> sigmoid(-5.65) = 0.00350519
        32'hC0B47AE1: sigmoid_out = 32'h3B680437; // -5.64 -> sigmoid(-5.64) = 0.00354029
        32'hC0B428F6: sigmoid_out = 32'h3B6A5705; // -5.63 -> sigmoid(-5.63) = 0.00357574
        32'hC0B3D70A: sigmoid_out = 32'h3B6CAFC3; // -5.62 -> sigmoid(-5.62) = 0.00361155
        32'hC0B3851F: sigmoid_out = 32'h3B6F0E80; // -5.61 -> sigmoid(-5.61) = 0.00364771
        32'hC0B33333: sigmoid_out = 32'h3B71734A; // -5.60 -> sigmoid(-5.60) = 0.00368424
        32'hC0B2E148: sigmoid_out = 32'h3B73DE31; // -5.59 -> sigmoid(-5.59) = 0.00372113
        32'hC0B28F5C: sigmoid_out = 32'h3B764F44; // -5.58 -> sigmoid(-5.58) = 0.00375839
        32'hC0B23D71: sigmoid_out = 32'h3B78C694; // -5.57 -> sigmoid(-5.57) = 0.00379602
        32'hC0B1EB85: sigmoid_out = 32'h3B7B442F; // -5.56 -> sigmoid(-5.56) = 0.00383402
        32'hC0B1999A: sigmoid_out = 32'h3B7DC826; // -5.55 -> sigmoid(-5.55) = 0.00387240
        32'hC0B147AE: sigmoid_out = 32'h3B802945; // -5.54 -> sigmoid(-5.54) = 0.00391117
        32'hC0B0F5C3: sigmoid_out = 32'h3B8171B4; // -5.53 -> sigmoid(-5.53) = 0.00395032
        32'hC0B0A3D7: sigmoid_out = 32'h3B82BD6A; // -5.52 -> sigmoid(-5.52) = 0.00398987
        32'hC0B051EC: sigmoid_out = 32'h3B840C6F; // -5.51 -> sigmoid(-5.51) = 0.00402980
        32'hC0B00000: sigmoid_out = 32'h3B855ECA; // -5.50 -> sigmoid(-5.50) = 0.00407014
        32'hC0AFAE14: sigmoid_out = 32'h3B86B485; // -5.49 -> sigmoid(-5.49) = 0.00411088
        32'hC0AF5C29: sigmoid_out = 32'h3B880DA8; // -5.48 -> sigmoid(-5.48) = 0.00415202
        32'hC0AF0A3D: sigmoid_out = 32'h3B896A3B; // -5.47 -> sigmoid(-5.47) = 0.00419357
        32'hC0AEB852: sigmoid_out = 32'h3B8ACA48; // -5.46 -> sigmoid(-5.46) = 0.00423554
        32'hC0AE6666: sigmoid_out = 32'h3B8C2DD7; // -5.45 -> sigmoid(-5.45) = 0.00427793
        32'hC0AE147B: sigmoid_out = 32'h3B8D94F1; // -5.44 -> sigmoid(-5.44) = 0.00432073
        32'hC0ADC28F: sigmoid_out = 32'h3B8EFF9E; // -5.43 -> sigmoid(-5.43) = 0.00436397
        32'hC0AD70A4: sigmoid_out = 32'h3B906DE9; // -5.42 -> sigmoid(-5.42) = 0.00440763
        32'hC0AD1EB8: sigmoid_out = 32'h3B91DFD9; // -5.41 -> sigmoid(-5.41) = 0.00445173
        32'hC0ACCCCD: sigmoid_out = 32'h3B935579; // -5.40 -> sigmoid(-5.40) = 0.00449627
        32'hC0AC7AE1: sigmoid_out = 32'h3B94CED2; // -5.39 -> sigmoid(-5.39) = 0.00454126
        32'hC0AC28F6: sigmoid_out = 32'h3B964BEC; // -5.38 -> sigmoid(-5.38) = 0.00458669
        32'hC0ABD70A: sigmoid_out = 32'h3B97CCD2; // -5.37 -> sigmoid(-5.37) = 0.00463257
        32'hC0AB851F: sigmoid_out = 32'h3B99518D; // -5.36 -> sigmoid(-5.36) = 0.00467891
        32'hC0AB3333: sigmoid_out = 32'h3B9ADA27; // -5.35 -> sigmoid(-5.35) = 0.00472571
        32'hC0AAE148: sigmoid_out = 32'h3B9C66A9; // -5.34 -> sigmoid(-5.34) = 0.00477298
        32'hC0AA8F5C: sigmoid_out = 32'h3B9DF71D; // -5.33 -> sigmoid(-5.33) = 0.00482072
        32'hC0AA3D71: sigmoid_out = 32'h3B9F8B8E; // -5.32 -> sigmoid(-5.32) = 0.00486893
        32'hC0A9EB85: sigmoid_out = 32'h3BA12406; // -5.31 -> sigmoid(-5.31) = 0.00491762
        32'hC0A9999A: sigmoid_out = 32'h3BA2C08D; // -5.30 -> sigmoid(-5.30) = 0.00496680
        32'hC0A947AE: sigmoid_out = 32'h3BA46130; // -5.29 -> sigmoid(-5.29) = 0.00501647
        32'hC0A8F5C3: sigmoid_out = 32'h3BA605F8; // -5.28 -> sigmoid(-5.28) = 0.00506663
        32'hC0A8A3D7: sigmoid_out = 32'h3BA7AEEF; // -5.27 -> sigmoid(-5.27) = 0.00511729
        32'hC0A851EC: sigmoid_out = 32'h3BA95C20; // -5.26 -> sigmoid(-5.26) = 0.00516845
        32'hC0A80000: sigmoid_out = 32'h3BAB0D97; // -5.25 -> sigmoid(-5.25) = 0.00522013
        32'hC0A7AE14: sigmoid_out = 32'h3BACC35C; // -5.24 -> sigmoid(-5.24) = 0.00527231
        32'hC0A75C29: sigmoid_out = 32'h3BAE7D7C; // -5.23 -> sigmoid(-5.23) = 0.00532502
        32'hC0A70A3D: sigmoid_out = 32'h3BB03C02; // -5.22 -> sigmoid(-5.22) = 0.00537825
        32'hC0A6B852: sigmoid_out = 32'h3BB1FEF8; // -5.21 -> sigmoid(-5.21) = 0.00543201
        32'hC0A66666: sigmoid_out = 32'h3BB3C669; // -5.20 -> sigmoid(-5.20) = 0.00548630
        32'hC0A6147B: sigmoid_out = 32'h3BB59261; // -5.19 -> sigmoid(-5.19) = 0.00554113
        32'hC0A5C28F: sigmoid_out = 32'h3BB762EC; // -5.18 -> sigmoid(-5.18) = 0.00559651
        32'hC0A570A4: sigmoid_out = 32'h3BB93814; // -5.17 -> sigmoid(-5.17) = 0.00565244
        32'hC0A51EB8: sigmoid_out = 32'h3BBB11E6; // -5.16 -> sigmoid(-5.16) = 0.00570892
        32'hC0A4CCCD: sigmoid_out = 32'h3BBCF06D; // -5.15 -> sigmoid(-5.15) = 0.00576597
        32'hC0A47AE1: sigmoid_out = 32'h3BBED3B4; // -5.14 -> sigmoid(-5.14) = 0.00582358
        32'hC0A428F6: sigmoid_out = 32'h3BC0BBC9; // -5.13 -> sigmoid(-5.13) = 0.00588176
        32'hC0A3D70A: sigmoid_out = 32'h3BC2A8B6; // -5.12 -> sigmoid(-5.12) = 0.00594052
        32'hC0A3851F: sigmoid_out = 32'h3BC49A89; // -5.11 -> sigmoid(-5.11) = 0.00599987
        32'hC0A33333: sigmoid_out = 32'h3BC6914D; // -5.10 -> sigmoid(-5.10) = 0.00605980
        32'hC0A2E148: sigmoid_out = 32'h3BC88D0E; // -5.09 -> sigmoid(-5.09) = 0.00612033
        32'hC0A28F5C: sigmoid_out = 32'h3BCA8DDA; // -5.08 -> sigmoid(-5.08) = 0.00618146
        32'hC0A23D71: sigmoid_out = 32'h3BCC93BD; // -5.07 -> sigmoid(-5.07) = 0.00624320
        32'hC0A1EB85: sigmoid_out = 32'h3BCE9EC4; // -5.06 -> sigmoid(-5.06) = 0.00630555
        32'hC0A1999A: sigmoid_out = 32'h3BD0AEFB; // -5.05 -> sigmoid(-5.05) = 0.00636852
        32'hC0A147AE: sigmoid_out = 32'h3BD2C470; // -5.04 -> sigmoid(-5.04) = 0.00643211
        32'hC0A0F5C3: sigmoid_out = 32'h3BD4DF2F; // -5.03 -> sigmoid(-5.03) = 0.00649633
        32'hC0A0A3D7: sigmoid_out = 32'h3BD6FF47; // -5.02 -> sigmoid(-5.02) = 0.00656119
        32'hC0A051EC: sigmoid_out = 32'h3BD924C4; // -5.01 -> sigmoid(-5.01) = 0.00662670
        32'hC0A00000: sigmoid_out = 32'h3BDB4FB4; // -5.00 -> sigmoid(-5.00) = 0.00669285
        32'hC09FAE14: sigmoid_out = 32'h3BDD8024; // -4.99 -> sigmoid(-4.99) = 0.00675966
        32'hC09F5C29: sigmoid_out = 32'h3BDFB623; // -4.98 -> sigmoid(-4.98) = 0.00682713
        32'hC09F0A3D: sigmoid_out = 32'h3BE1F1BE; // -4.97 -> sigmoid(-4.97) = 0.00689527
        32'hC09EB852: sigmoid_out = 32'h3BE43304; // -4.96 -> sigmoid(-4.96) = 0.00696409
        32'hC09E6666: sigmoid_out = 32'h3BE67A01; // -4.95 -> sigmoid(-4.95) = 0.00703359
        32'hC09E147B: sigmoid_out = 32'h3BE8C6C6; // -4.94 -> sigmoid(-4.94) = 0.00710377
        32'hC09DC28F: sigmoid_out = 32'h3BEB1960; // -4.93 -> sigmoid(-4.93) = 0.00717466
        32'hC09D70A4: sigmoid_out = 32'h3BED71DD; // -4.92 -> sigmoid(-4.92) = 0.00724624
        32'hC09D1EB8: sigmoid_out = 32'h3BEFD04D; // -4.91 -> sigmoid(-4.91) = 0.00731853
        32'hC09CCCCD: sigmoid_out = 32'h3BF234BE; // -4.90 -> sigmoid(-4.90) = 0.00739154
        32'hC09C7AE1: sigmoid_out = 32'h3BF49F40; // -4.89 -> sigmoid(-4.89) = 0.00746527
        32'hC09C28F6: sigmoid_out = 32'h3BF70FE1; // -4.88 -> sigmoid(-4.88) = 0.00753973
        32'hC09BD70A: sigmoid_out = 32'h3BF986B0; // -4.87 -> sigmoid(-4.87) = 0.00761493
        32'hC09B851F: sigmoid_out = 32'h3BFC03BE; // -4.86 -> sigmoid(-4.86) = 0.00769088
        32'hC09B3333: sigmoid_out = 32'h3BFE871A; // -4.85 -> sigmoid(-4.85) = 0.00776757
        32'hC09AE148: sigmoid_out = 32'h3C008869; // -4.84 -> sigmoid(-4.84) = 0.00784502
        32'hC09A8F5C: sigmoid_out = 32'h3C01D07C; // -4.83 -> sigmoid(-4.83) = 0.00792324
        32'hC09A3D71: sigmoid_out = 32'h3C031BCE; // -4.82 -> sigmoid(-4.82) = 0.00800223
        32'hC099EB85: sigmoid_out = 32'h3C046A67; // -4.81 -> sigmoid(-4.81) = 0.00808201
        32'hC099999A: sigmoid_out = 32'h3C05BC4E; // -4.80 -> sigmoid(-4.80) = 0.00816257
        32'hC09947AE: sigmoid_out = 32'h3C07118D; // -4.79 -> sigmoid(-4.79) = 0.00824393
        32'hC098F5C3: sigmoid_out = 32'h3C086A2A; // -4.78 -> sigmoid(-4.78) = 0.00832609
        32'hC098A3D7: sigmoid_out = 32'h3C09C630; // -4.77 -> sigmoid(-4.77) = 0.00840907
        32'hC09851EC: sigmoid_out = 32'h3C0B25A6; // -4.76 -> sigmoid(-4.76) = 0.00849286
        32'hC0980000: sigmoid_out = 32'h3C0C8895; // -4.75 -> sigmoid(-4.75) = 0.00857749
        32'hC097AE14: sigmoid_out = 32'h3C0DEF05; // -4.74 -> sigmoid(-4.74) = 0.00866294
        32'hC0975C29: sigmoid_out = 32'h3C0F58FF; // -4.73 -> sigmoid(-4.73) = 0.00874925
        32'hC0970A3D: sigmoid_out = 32'h3C10C68D; // -4.72 -> sigmoid(-4.72) = 0.00883640
        32'hC096B852: sigmoid_out = 32'h3C1237B6; // -4.71 -> sigmoid(-4.71) = 0.00892442
        32'hC0966666: sigmoid_out = 32'h3C13AC84; // -4.70 -> sigmoid(-4.70) = 0.00901330
        32'hC096147B: sigmoid_out = 32'h3C1524FF; // -4.69 -> sigmoid(-4.69) = 0.00910306
        32'hC095C28F: sigmoid_out = 32'h3C16A132; // -4.68 -> sigmoid(-4.68) = 0.00919371
        32'hC09570A4: sigmoid_out = 32'h3C182125; // -4.67 -> sigmoid(-4.67) = 0.00928525
        32'hC0951EB8: sigmoid_out = 32'h3C19A4E1; // -4.66 -> sigmoid(-4.66) = 0.00937769
        32'hC094CCCD: sigmoid_out = 32'h3C1B2C70; // -4.65 -> sigmoid(-4.65) = 0.00947104
        32'hC0947AE1: sigmoid_out = 32'h3C1CB7DB; // -4.64 -> sigmoid(-4.64) = 0.00956532
        32'hC09428F6: sigmoid_out = 32'h3C1E472C; // -4.63 -> sigmoid(-4.63) = 0.00966052
        32'hC093D70A: sigmoid_out = 32'h3C1FDA6C; // -4.62 -> sigmoid(-4.62) = 0.00975667
        32'hC093851F: sigmoid_out = 32'h3C2171A5; // -4.61 -> sigmoid(-4.61) = 0.00985376
        32'hC0933333: sigmoid_out = 32'h3C230CE2; // -4.60 -> sigmoid(-4.60) = 0.00995180
        32'hC092E148: sigmoid_out = 32'h3C24AC2B; // -4.59 -> sigmoid(-4.59) = 0.01005081
        32'hC0928F5C: sigmoid_out = 32'h3C264F8B; // -4.58 -> sigmoid(-4.58) = 0.01015080
        32'hC0923D71: sigmoid_out = 32'h3C27F70D; // -4.57 -> sigmoid(-4.57) = 0.01025177
        32'hC091EB85: sigmoid_out = 32'h3C29A2B9; // -4.56 -> sigmoid(-4.56) = 0.01035374
        32'hC091999A: sigmoid_out = 32'h3C2B529B; // -4.55 -> sigmoid(-4.55) = 0.01045671
        32'hC09147AE: sigmoid_out = 32'h3C2D06BC; // -4.54 -> sigmoid(-4.54) = 0.01056069
        32'hC090F5C3: sigmoid_out = 32'h3C2EBF28; // -4.53 -> sigmoid(-4.53) = 0.01066569
        32'hC090A3D7: sigmoid_out = 32'h3C307BE9; // -4.52 -> sigmoid(-4.52) = 0.01077173
        32'hC09051EC: sigmoid_out = 32'h3C323D09; // -4.51 -> sigmoid(-4.51) = 0.01087881
        32'hC0900000: sigmoid_out = 32'h3C340294; // -4.50 -> sigmoid(-4.50) = 0.01098694
        32'hC08FAE14: sigmoid_out = 32'h3C35CC93; // -4.49 -> sigmoid(-4.49) = 0.01109614
        32'hC08F5C29: sigmoid_out = 32'h3C379B13; // -4.48 -> sigmoid(-4.48) = 0.01120641
        32'hC08F0A3D: sigmoid_out = 32'h3C396E1E; // -4.47 -> sigmoid(-4.47) = 0.01131776
        32'hC08EB852: sigmoid_out = 32'h3C3B45BF; // -4.46 -> sigmoid(-4.46) = 0.01143020
        32'hC08E6666: sigmoid_out = 32'h3C3D2202; // -4.45 -> sigmoid(-4.45) = 0.01154375
        32'hC08E147B: sigmoid_out = 32'h3C3F02F1; // -4.44 -> sigmoid(-4.44) = 0.01165842
        32'hC08DC28F: sigmoid_out = 32'h3C40E899; // -4.43 -> sigmoid(-4.43) = 0.01177421
        32'hC08D70A4: sigmoid_out = 32'h3C42D305; // -4.42 -> sigmoid(-4.42) = 0.01189113
        32'hC08D1EB8: sigmoid_out = 32'h3C44C241; // -4.41 -> sigmoid(-4.41) = 0.01200920
        32'hC08CCCCD: sigmoid_out = 32'h3C46B658; // -4.40 -> sigmoid(-4.40) = 0.01212843
        32'hC08C7AE1: sigmoid_out = 32'h3C48AF56; // -4.39 -> sigmoid(-4.39) = 0.01224883
        32'hC08C28F6: sigmoid_out = 32'h3C4AAD48; // -4.38 -> sigmoid(-4.38) = 0.01237041
        32'hC08BD70A: sigmoid_out = 32'h3C4CB039; // -4.37 -> sigmoid(-4.37) = 0.01249319
        32'hC08B851F: sigmoid_out = 32'h3C4EB835; // -4.36 -> sigmoid(-4.36) = 0.01261716
        32'hC08B3333: sigmoid_out = 32'h3C50C54A; // -4.35 -> sigmoid(-4.35) = 0.01274235
        32'hC08AE148: sigmoid_out = 32'h3C52D782; // -4.34 -> sigmoid(-4.34) = 0.01286876
        32'hC08A8F5C: sigmoid_out = 32'h3C54EEEC; // -4.33 -> sigmoid(-4.33) = 0.01299642
        32'hC08A3D71: sigmoid_out = 32'h3C570B93; // -4.32 -> sigmoid(-4.32) = 0.01312532
        32'hC089EB85: sigmoid_out = 32'h3C592D85; // -4.31 -> sigmoid(-4.31) = 0.01325548
        32'hC089999A: sigmoid_out = 32'h3C5B54CE; // -4.30 -> sigmoid(-4.30) = 0.01338692
        32'hC08947AE: sigmoid_out = 32'h3C5D817B; // -4.29 -> sigmoid(-4.29) = 0.01351964
        32'hC088F5C3: sigmoid_out = 32'h3C5FB399; // -4.28 -> sigmoid(-4.28) = 0.01365366
        32'hC088A3D7: sigmoid_out = 32'h3C61EB36; // -4.27 -> sigmoid(-4.27) = 0.01378899
        32'hC08851EC: sigmoid_out = 32'h3C64285E; // -4.26 -> sigmoid(-4.26) = 0.01392564
        32'hC0880000: sigmoid_out = 32'h3C666B21; // -4.25 -> sigmoid(-4.25) = 0.01406363
        32'hC087AE14: sigmoid_out = 32'h3C68B38A; // -4.24 -> sigmoid(-4.24) = 0.01420296
        32'hC0875C29: sigmoid_out = 32'h3C6B01A7; // -4.23 -> sigmoid(-4.23) = 0.01434366
        32'hC0870A3D: sigmoid_out = 32'h3C6D5588; // -4.22 -> sigmoid(-4.22) = 0.01448572
        32'hC086B852: sigmoid_out = 32'h3C6FAF38; // -4.21 -> sigmoid(-4.21) = 0.01462918
        32'hC0866666: sigmoid_out = 32'h3C720EC8; // -4.20 -> sigmoid(-4.20) = 0.01477403
        32'hC086147B: sigmoid_out = 32'h3C747444; // -4.19 -> sigmoid(-4.19) = 0.01492030
        32'hC085C28F: sigmoid_out = 32'h3C76DFBB; // -4.18 -> sigmoid(-4.18) = 0.01506799
        32'hC08570A4: sigmoid_out = 32'h3C79513B; // -4.17 -> sigmoid(-4.17) = 0.01521712
        32'hC0851EB8: sigmoid_out = 32'h3C7BC8D4; // -4.16 -> sigmoid(-4.16) = 0.01536771
        32'hC084CCCD: sigmoid_out = 32'h3C7E4694; // -4.15 -> sigmoid(-4.15) = 0.01551976
        32'hC0847AE1: sigmoid_out = 32'h3C806544; // -4.14 -> sigmoid(-4.14) = 0.01567329
        32'hC08428F6: sigmoid_out = 32'h3C81AA61; // -4.13 -> sigmoid(-4.13) = 0.01582831
        32'hC083D70A: sigmoid_out = 32'h3C82F2A8; // -4.12 -> sigmoid(-4.12) = 0.01598485
        32'hC083851F: sigmoid_out = 32'h3C843E20; // -4.11 -> sigmoid(-4.11) = 0.01614291
        32'hC0833333: sigmoid_out = 32'h3C858CD2; // -4.10 -> sigmoid(-4.10) = 0.01630250
        32'hC082E148: sigmoid_out = 32'h3C86DEC4; // -4.09 -> sigmoid(-4.09) = 0.01646364
        32'hC0828F5C: sigmoid_out = 32'h3C8833FF; // -4.08 -> sigmoid(-4.08) = 0.01662636
        32'hC0823D71: sigmoid_out = 32'h3C898C8B; // -4.07 -> sigmoid(-4.07) = 0.01679065
        32'hC081EB85: sigmoid_out = 32'h3C8AE86F; // -4.06 -> sigmoid(-4.06) = 0.01695654
        32'hC081999A: sigmoid_out = 32'h3C8C47B3; // -4.05 -> sigmoid(-4.05) = 0.01712403
        32'hC08147AE: sigmoid_out = 32'h3C8DAA61; // -4.04 -> sigmoid(-4.04) = 0.01729316
        32'hC080F5C3: sigmoid_out = 32'h3C8F107F; // -4.03 -> sigmoid(-4.03) = 0.01746392
        32'hC080A3D7: sigmoid_out = 32'h3C907A16; // -4.02 -> sigmoid(-4.02) = 0.01763634
        32'hC08051EC: sigmoid_out = 32'h3C91E72F; // -4.01 -> sigmoid(-4.01) = 0.01781043
        32'hC0800000: sigmoid_out = 32'h3C9357D1; // -4.00 -> sigmoid(-4.00) = 0.01798621
        32'hC07F5C29: sigmoid_out = 32'h3C94CC05; // -3.99 -> sigmoid(-3.99) = 0.01816369
        32'hC07EB852: sigmoid_out = 32'h3C9643D4; // -3.98 -> sigmoid(-3.98) = 0.01834289
        32'hC07E147B: sigmoid_out = 32'h3C97BF47; // -3.97 -> sigmoid(-3.97) = 0.01852382
        32'hC07D70A4: sigmoid_out = 32'h3C993E65; // -3.96 -> sigmoid(-3.96) = 0.01870651
        32'hC07CCCCD: sigmoid_out = 32'h3C9AC138; // -3.95 -> sigmoid(-3.95) = 0.01889096
        32'hC07C28F6: sigmoid_out = 32'h3C9C47C8; // -3.94 -> sigmoid(-3.94) = 0.01907720
        32'hC07B851F: sigmoid_out = 32'h3C9DD21F; // -3.93 -> sigmoid(-3.93) = 0.01926523
        32'hC07AE148: sigmoid_out = 32'h3C9F6045; // -3.92 -> sigmoid(-3.92) = 0.01945508
        32'hC07A3D71: sigmoid_out = 32'h3CA0F243; // -3.91 -> sigmoid(-3.91) = 0.01964677
        32'hC079999A: sigmoid_out = 32'h3CA28823; // -3.90 -> sigmoid(-3.90) = 0.01984031
        32'hC078F5C3: sigmoid_out = 32'h3CA421ED; // -3.89 -> sigmoid(-3.89) = 0.02003571
        32'hC07851EC: sigmoid_out = 32'h3CA5BFAC; // -3.88 -> sigmoid(-3.88) = 0.02023300
        32'hC077AE14: sigmoid_out = 32'h3CA76167; // -3.87 -> sigmoid(-3.87) = 0.02043219
        32'hC0770A3D: sigmoid_out = 32'h3CA90729; // -3.86 -> sigmoid(-3.86) = 0.02063330
        32'hC0766666: sigmoid_out = 32'h3CAAB0FB; // -3.85 -> sigmoid(-3.85) = 0.02083634
        32'hC075C28F: sigmoid_out = 32'h3CAC5EE7; // -3.84 -> sigmoid(-3.84) = 0.02104135
        32'hC0751EB8: sigmoid_out = 32'h3CAE10F6; // -3.83 -> sigmoid(-3.83) = 0.02124832
        32'hC0747AE1: sigmoid_out = 32'h3CAFC733; // -3.82 -> sigmoid(-3.82) = 0.02145729
        32'hC073D70A: sigmoid_out = 32'h3CB181A6; // -3.81 -> sigmoid(-3.81) = 0.02166827
        32'hC0733333: sigmoid_out = 32'h3CB3405A; // -3.80 -> sigmoid(-3.80) = 0.02188127
        32'hC0728F5C: sigmoid_out = 32'h3CB50359; // -3.79 -> sigmoid(-3.79) = 0.02209632
        32'hC071EB85: sigmoid_out = 32'h3CB6CAAC; // -3.78 -> sigmoid(-3.78) = 0.02231344
        32'hC07147AE: sigmoid_out = 32'h3CB8965F; // -3.77 -> sigmoid(-3.77) = 0.02253264
        32'hC070A3D7: sigmoid_out = 32'h3CBA667A; // -3.76 -> sigmoid(-3.76) = 0.02275394
        32'hC0700000: sigmoid_out = 32'h3CBC3B0A; // -3.75 -> sigmoid(-3.75) = 0.02297737
        32'hC06F5C29: sigmoid_out = 32'h3CBE1417; // -3.74 -> sigmoid(-3.74) = 0.02320294
        32'hC06EB852: sigmoid_out = 32'h3CBFF1AC; // -3.73 -> sigmoid(-3.73) = 0.02343067
        32'hC06E147B: sigmoid_out = 32'h3CC1D3D4; // -3.72 -> sigmoid(-3.72) = 0.02366058
        32'hC06D70A4: sigmoid_out = 32'h3CC3BA9A; // -3.71 -> sigmoid(-3.71) = 0.02389269
        32'hC06CCCCD: sigmoid_out = 32'h3CC5A608; // -3.70 -> sigmoid(-3.70) = 0.02412702
        32'hC06C28F6: sigmoid_out = 32'h3CC79629; // -3.69 -> sigmoid(-3.69) = 0.02436359
        32'hC06B851F: sigmoid_out = 32'h3CC98B08; // -3.68 -> sigmoid(-3.68) = 0.02460243
        32'hC06AE148: sigmoid_out = 32'h3CCB84B0; // -3.67 -> sigmoid(-3.67) = 0.02484354
        32'hC06A3D71: sigmoid_out = 32'h3CCD832C; // -3.66 -> sigmoid(-3.66) = 0.02508696
        32'hC069999A: sigmoid_out = 32'h3CCF8687; // -3.65 -> sigmoid(-3.65) = 0.02533270
        32'hC068F5C3: sigmoid_out = 32'h3CD18ECD; // -3.64 -> sigmoid(-3.64) = 0.02558079
        32'hC06851EC: sigmoid_out = 32'h3CD39C09; // -3.63 -> sigmoid(-3.63) = 0.02583124
        32'hC067AE14: sigmoid_out = 32'h3CD5AE45; // -3.62 -> sigmoid(-3.62) = 0.02608408
        32'hC0670A3D: sigmoid_out = 32'h3CD7C58F; // -3.61 -> sigmoid(-3.61) = 0.02633932
        32'hC0666666: sigmoid_out = 32'h3CD9E1F0; // -3.60 -> sigmoid(-3.60) = 0.02659699
        32'hC065C28F: sigmoid_out = 32'h3CDC0376; // -3.59 -> sigmoid(-3.59) = 0.02685712
        32'hC0651EB8: sigmoid_out = 32'h3CDE2A2B; // -3.58 -> sigmoid(-3.58) = 0.02711972
        32'hC0647AE1: sigmoid_out = 32'h3CE0561C; // -3.57 -> sigmoid(-3.57) = 0.02738481
        32'hC063D70A: sigmoid_out = 32'h3CE28755; // -3.56 -> sigmoid(-3.56) = 0.02765242
        32'hC0633333: sigmoid_out = 32'h3CE4BDE2; // -3.55 -> sigmoid(-3.55) = 0.02792257
        32'hC0628F5C: sigmoid_out = 32'h3CE6F9CE; // -3.54 -> sigmoid(-3.54) = 0.02819529
        32'hC061EB85: sigmoid_out = 32'h3CE93B26; // -3.53 -> sigmoid(-3.53) = 0.02847059
        32'hC06147AE: sigmoid_out = 32'h3CEB81F7; // -3.52 -> sigmoid(-3.52) = 0.02874850
        32'hC060A3D7: sigmoid_out = 32'h3CEDCE4D; // -3.51 -> sigmoid(-3.51) = 0.02902904
        32'hC0600000: sigmoid_out = 32'h3CF02034; // -3.50 -> sigmoid(-3.50) = 0.02931223
        32'hC05F5C29: sigmoid_out = 32'h3CF277B9; // -3.49 -> sigmoid(-3.49) = 0.02959810
        32'hC05EB852: sigmoid_out = 32'h3CF4D4E9; // -3.48 -> sigmoid(-3.48) = 0.02988668
        32'hC05E147B: sigmoid_out = 32'h3CF737D0; // -3.47 -> sigmoid(-3.47) = 0.03017798
        32'hC05D70A4: sigmoid_out = 32'h3CF9A07C; // -3.46 -> sigmoid(-3.46) = 0.03047203
        32'hC05CCCCD: sigmoid_out = 32'h3CFC0EFA; // -3.45 -> sigmoid(-3.45) = 0.03076886
        32'hC05C28F6: sigmoid_out = 32'h3CFE8355; // -3.44 -> sigmoid(-3.44) = 0.03106848
        32'hC05B851F: sigmoid_out = 32'h3D007ECF; // -3.43 -> sigmoid(-3.43) = 0.03137093
        32'hC05AE148: sigmoid_out = 32'h3D01BEEF; // -3.42 -> sigmoid(-3.42) = 0.03167623
        32'hC05A3D71: sigmoid_out = 32'h3D030212; // -3.41 -> sigmoid(-3.41) = 0.03198440
        32'hC059999A: sigmoid_out = 32'h3D044840; // -3.40 -> sigmoid(-3.40) = 0.03229546
        32'hC058F5C3: sigmoid_out = 32'h3D05917E; // -3.39 -> sigmoid(-3.39) = 0.03260946
        32'hC05851EC: sigmoid_out = 32'h3D06DDD4; // -3.38 -> sigmoid(-3.38) = 0.03292639
        32'hC057AE14: sigmoid_out = 32'h3D082D48; // -3.37 -> sigmoid(-3.37) = 0.03324631
        32'hC0570A3D: sigmoid_out = 32'h3D097FE2; // -3.36 -> sigmoid(-3.36) = 0.03356922
        32'hC0566666: sigmoid_out = 32'h3D0AD5A8; // -3.35 -> sigmoid(-3.35) = 0.03389516
        32'hC055C28F: sigmoid_out = 32'h3D0C2EA1; // -3.34 -> sigmoid(-3.34) = 0.03422416
        32'hC0551EB8: sigmoid_out = 32'h3D0D8AD5; // -3.33 -> sigmoid(-3.33) = 0.03455623
        32'hC0547AE1: sigmoid_out = 32'h3D0EEA4B; // -3.32 -> sigmoid(-3.32) = 0.03489141
        32'hC053D70A: sigmoid_out = 32'h3D104D0A; // -3.31 -> sigmoid(-3.31) = 0.03522972
        32'hC0533333: sigmoid_out = 32'h3D11B318; // -3.30 -> sigmoid(-3.30) = 0.03557119
        32'hC0528F5C: sigmoid_out = 32'h3D131C7E; // -3.29 -> sigmoid(-3.29) = 0.03591585
        32'hC051EB85: sigmoid_out = 32'h3D148943; // -3.28 -> sigmoid(-3.28) = 0.03626372
        32'hC05147AE: sigmoid_out = 32'h3D15F96E; // -3.27 -> sigmoid(-3.27) = 0.03661483
        32'hC050A3D7: sigmoid_out = 32'h3D176D07; // -3.26 -> sigmoid(-3.26) = 0.03696921
        32'hC0500000: sigmoid_out = 32'h3D18E414; // -3.25 -> sigmoid(-3.25) = 0.03732689
        32'hC04F5C29: sigmoid_out = 32'h3D1A5E9E; // -3.24 -> sigmoid(-3.24) = 0.03768789
        32'hC04EB852: sigmoid_out = 32'h3D1BDCAC; // -3.23 -> sigmoid(-3.23) = 0.03805225
        32'hC04E147B: sigmoid_out = 32'h3D1D5E46; // -3.22 -> sigmoid(-3.22) = 0.03841999
        32'hC04D70A4: sigmoid_out = 32'h3D1EE374; // -3.21 -> sigmoid(-3.21) = 0.03879113
        32'hC04CCCCD: sigmoid_out = 32'h3D206C3D; // -3.20 -> sigmoid(-3.20) = 0.03916572
        32'hC04C28F6: sigmoid_out = 32'h3D21F8A8; // -3.19 -> sigmoid(-3.19) = 0.03954378
        32'hC04B851F: sigmoid_out = 32'h3D2388BF; // -3.18 -> sigmoid(-3.18) = 0.03992533
        32'hC04AE148: sigmoid_out = 32'h3D251C89; // -3.17 -> sigmoid(-3.17) = 0.04031042
        32'hC04A3D71: sigmoid_out = 32'h3D26B40D; // -3.16 -> sigmoid(-3.16) = 0.04069905
        32'hC049999A: sigmoid_out = 32'h3D284F54; // -3.15 -> sigmoid(-3.15) = 0.04109128
        32'hC048F5C3: sigmoid_out = 32'h3D29EE66; // -3.14 -> sigmoid(-3.14) = 0.04148712
        32'hC04851EC: sigmoid_out = 32'h3D2B914A; // -3.13 -> sigmoid(-3.13) = 0.04188661
        32'hC047AE14: sigmoid_out = 32'h3D2D380A; // -3.12 -> sigmoid(-3.12) = 0.04228977
        32'hC0470A3D: sigmoid_out = 32'h3D2EE2AD; // -3.11 -> sigmoid(-3.11) = 0.04269664
        32'hC0466666: sigmoid_out = 32'h3D30913C; // -3.10 -> sigmoid(-3.10) = 0.04310725
        32'hC045C28F: sigmoid_out = 32'h3D3243BE; // -3.09 -> sigmoid(-3.09) = 0.04352163
        32'hC0451EB8: sigmoid_out = 32'h3D33FA3C; // -3.08 -> sigmoid(-3.08) = 0.04393982
        32'hC0447AE1: sigmoid_out = 32'h3D35B4BF; // -3.07 -> sigmoid(-3.07) = 0.04436183
        32'hC043D70A: sigmoid_out = 32'h3D37734F; // -3.06 -> sigmoid(-3.06) = 0.04478770
        32'hC0433333: sigmoid_out = 32'h3D3935F5; // -3.05 -> sigmoid(-3.05) = 0.04521747
        32'hC0428F5C: sigmoid_out = 32'h3D3AFCB9; // -3.04 -> sigmoid(-3.04) = 0.04565117
        32'hC041EB85: sigmoid_out = 32'h3D3CC7A3; // -3.03 -> sigmoid(-3.03) = 0.04608883
        32'hC04147AE: sigmoid_out = 32'h3D3E96BD; // -3.02 -> sigmoid(-3.02) = 0.04653047
        32'hC040A3D7: sigmoid_out = 32'h3D406A0F; // -3.01 -> sigmoid(-3.01) = 0.04697615
        32'hC0400000: sigmoid_out = 32'h3D4241A2; // -3.00 -> sigmoid(-3.00) = 0.04742587
        32'hC03F5C29: sigmoid_out = 32'h3D441D7E; // -2.99 -> sigmoid(-2.99) = 0.04787969
        32'hC03EB852: sigmoid_out = 32'h3D45FDAD; // -2.98 -> sigmoid(-2.98) = 0.04833763
        32'hC03E147B: sigmoid_out = 32'h3D47E238; // -2.97 -> sigmoid(-2.97) = 0.04879972
        32'hC03D70A4: sigmoid_out = 32'h3D49CB27; // -2.96 -> sigmoid(-2.96) = 0.04926601
        32'hC03CCCCD: sigmoid_out = 32'h3D4BB883; // -2.95 -> sigmoid(-2.95) = 0.04973651
        32'hC03C28F6: sigmoid_out = 32'h3D4DAA56; // -2.94 -> sigmoid(-2.94) = 0.05021127
        32'hC03B851F: sigmoid_out = 32'h3D4FA0A8; // -2.93 -> sigmoid(-2.93) = 0.05069032
        32'hC03AE148: sigmoid_out = 32'h3D519B84; // -2.92 -> sigmoid(-2.92) = 0.05117370
        32'hC03A3D71: sigmoid_out = 32'h3D539AF1; // -2.91 -> sigmoid(-2.91) = 0.05166144
        32'hC039999A: sigmoid_out = 32'h3D559EF9; // -2.90 -> sigmoid(-2.90) = 0.05215356
        32'hC038F5C3: sigmoid_out = 32'h3D57A7A7; // -2.89 -> sigmoid(-2.89) = 0.05265012
        32'hC03851EC: sigmoid_out = 32'h3D59B502; // -2.88 -> sigmoid(-2.88) = 0.05315114
        32'hC037AE14: sigmoid_out = 32'h3D5BC714; // -2.87 -> sigmoid(-2.87) = 0.05365665
        32'hC0370A3D: sigmoid_out = 32'h3D5DDDE7; // -2.86 -> sigmoid(-2.86) = 0.05416670
        32'hC0366666: sigmoid_out = 32'h3D5FF984; // -2.85 -> sigmoid(-2.85) = 0.05468132
        32'hC035C28F: sigmoid_out = 32'h3D6219F6; // -2.84 -> sigmoid(-2.84) = 0.05520054
        32'hC0351EB8: sigmoid_out = 32'h3D643F44; // -2.83 -> sigmoid(-2.83) = 0.05572440
        32'hC0347AE1: sigmoid_out = 32'h3D66697A; // -2.82 -> sigmoid(-2.82) = 0.05625293
        32'hC033D70A: sigmoid_out = 32'h3D6898A0; // -2.81 -> sigmoid(-2.81) = 0.05678618
        32'hC0333333: sigmoid_out = 32'h3D6ACCC1; // -2.80 -> sigmoid(-2.80) = 0.05732418
        32'hC0328F5C: sigmoid_out = 32'h3D6D05E7; // -2.79 -> sigmoid(-2.79) = 0.05786696
        32'hC031EB85: sigmoid_out = 32'h3D6F441A; // -2.78 -> sigmoid(-2.78) = 0.05841456
        32'hC03147AE: sigmoid_out = 32'h3D718765; // -2.77 -> sigmoid(-2.77) = 0.05896701
        32'hC030A3D7: sigmoid_out = 32'h3D73CFD2; // -2.76 -> sigmoid(-2.76) = 0.05952437
        32'hC0300000: sigmoid_out = 32'h3D761D6B; // -2.75 -> sigmoid(-2.75) = 0.06008665
        32'hC02F5C29: sigmoid_out = 32'h3D78703A; // -2.74 -> sigmoid(-2.74) = 0.06065390
        32'hC02EB852: sigmoid_out = 32'h3D7AC849; // -2.73 -> sigmoid(-2.73) = 0.06122616
        32'hC02E147B: sigmoid_out = 32'h3D7D25A2; // -2.72 -> sigmoid(-2.72) = 0.06180347
        32'hC02D70A4: sigmoid_out = 32'h3D7F884E; // -2.71 -> sigmoid(-2.71) = 0.06238585
        32'hC02CCCCD: sigmoid_out = 32'h3D80F82D; // -2.70 -> sigmoid(-2.70) = 0.06297336
        32'hC02C28F6: sigmoid_out = 32'h3D822EE7; // -2.69 -> sigmoid(-2.69) = 0.06356602
        32'hC02B851F: sigmoid_out = 32'h3D83685A; // -2.68 -> sigmoid(-2.68) = 0.06416388
        32'hC02AE148: sigmoid_out = 32'h3D84A48B; // -2.67 -> sigmoid(-2.67) = 0.06476697
        32'hC02A3D71: sigmoid_out = 32'h3D85E381; // -2.66 -> sigmoid(-2.66) = 0.06537533
        32'hC029999A: sigmoid_out = 32'h3D87253F; // -2.65 -> sigmoid(-2.65) = 0.06598901
        32'hC028F5C3: sigmoid_out = 32'h3D8869CB; // -2.64 -> sigmoid(-2.64) = 0.06660804
        32'hC02851EC: sigmoid_out = 32'h3D89B12B; // -2.63 -> sigmoid(-2.63) = 0.06723245
        32'hC027AE14: sigmoid_out = 32'h3D8AFB63; // -2.62 -> sigmoid(-2.62) = 0.06786229
        32'hC0270A3D: sigmoid_out = 32'h3D8C4879; // -2.61 -> sigmoid(-2.61) = 0.06849760
        32'hC0266666: sigmoid_out = 32'h3D8D9872; // -2.60 -> sigmoid(-2.60) = 0.06913842
        32'hC025C28F: sigmoid_out = 32'h3D8EEB53; // -2.59 -> sigmoid(-2.59) = 0.06978478
        32'hC0251EB8: sigmoid_out = 32'h3D904122; // -2.58 -> sigmoid(-2.58) = 0.07043673
        32'hC0247AE1: sigmoid_out = 32'h3D9199E4; // -2.57 -> sigmoid(-2.57) = 0.07109430
        32'hC023D70A: sigmoid_out = 32'h3D92F59E; // -2.56 -> sigmoid(-2.56) = 0.07175754
        32'hC0233333: sigmoid_out = 32'h3D945456; // -2.55 -> sigmoid(-2.55) = 0.07242649
        32'hC0228F5C: sigmoid_out = 32'h3D95B611; // -2.54 -> sigmoid(-2.54) = 0.07310117
        32'hC021EB85: sigmoid_out = 32'h3D971AD5; // -2.53 -> sigmoid(-2.53) = 0.07378165
        32'hC02147AE: sigmoid_out = 32'h3D9882A6; // -2.52 -> sigmoid(-2.52) = 0.07446795
        32'hC020A3D7: sigmoid_out = 32'h3D99ED8B; // -2.51 -> sigmoid(-2.51) = 0.07516011
        32'hC0200000: sigmoid_out = 32'h3D9B5B89; // -2.50 -> sigmoid(-2.50) = 0.07585818
        32'hC01F5C29: sigmoid_out = 32'h3D9CCCA4; // -2.49 -> sigmoid(-2.49) = 0.07656220
        32'hC01EB852: sigmoid_out = 32'h3D9E40E3; // -2.48 -> sigmoid(-2.48) = 0.07727220
        32'hC01E147B: sigmoid_out = 32'h3D9FB84C; // -2.47 -> sigmoid(-2.47) = 0.07798824
        32'hC01D70A4: sigmoid_out = 32'h3DA132E3; // -2.46 -> sigmoid(-2.46) = 0.07871034
        32'hC01CCCCD: sigmoid_out = 32'h3DA2B0AE; // -2.45 -> sigmoid(-2.45) = 0.07943855
        32'hC01C28F6: sigmoid_out = 32'h3DA431B2; // -2.44 -> sigmoid(-2.44) = 0.08017291
        32'hC01B851F: sigmoid_out = 32'h3DA5B5F6; // -2.43 -> sigmoid(-2.43) = 0.08091347
        32'hC01AE148: sigmoid_out = 32'h3DA73D7E; // -2.42 -> sigmoid(-2.42) = 0.08166026
        32'hC01A3D71: sigmoid_out = 32'h3DA8C850; // -2.41 -> sigmoid(-2.41) = 0.08241332
        32'hC019999A: sigmoid_out = 32'h3DAA5672; // -2.40 -> sigmoid(-2.40) = 0.08317270
        32'hC018F5C3: sigmoid_out = 32'h3DABE7EA; // -2.39 -> sigmoid(-2.39) = 0.08393843
        32'hC01851EC: sigmoid_out = 32'h3DAD7CBC; // -2.38 -> sigmoid(-2.38) = 0.08471057
        32'hC017AE14: sigmoid_out = 32'h3DAF14EE; // -2.37 -> sigmoid(-2.37) = 0.08548914
        32'hC0170A3D: sigmoid_out = 32'h3DB0B086; // -2.36 -> sigmoid(-2.36) = 0.08627419
        32'hC0166666: sigmoid_out = 32'h3DB24F8A; // -2.35 -> sigmoid(-2.35) = 0.08706577
        32'hC015C28F: sigmoid_out = 32'h3DB3F1FF; // -2.34 -> sigmoid(-2.34) = 0.08786391
        32'hC0151EB8: sigmoid_out = 32'h3DB597EB; // -2.33 -> sigmoid(-2.33) = 0.08866866
        32'hC0147AE1: sigmoid_out = 32'h3DB74152; // -2.32 -> sigmoid(-2.32) = 0.08948006
        32'hC013D70A: sigmoid_out = 32'h3DB8EE3C; // -2.31 -> sigmoid(-2.31) = 0.09029814
        32'hC0133333: sigmoid_out = 32'h3DBA9EAD; // -2.30 -> sigmoid(-2.30) = 0.09112296
        32'hC0128F5C: sigmoid_out = 32'h3DBC52AB; // -2.29 -> sigmoid(-2.29) = 0.09195455
        32'hC011EB85: sigmoid_out = 32'h3DBE0A3B; // -2.28 -> sigmoid(-2.28) = 0.09279295
        32'hC01147AE: sigmoid_out = 32'h3DBFC564; // -2.27 -> sigmoid(-2.27) = 0.09363821
        32'hC010A3D7: sigmoid_out = 32'h3DC1842B; // -2.26 -> sigmoid(-2.26) = 0.09449037
        32'hC0100000: sigmoid_out = 32'h3DC34695; // -2.25 -> sigmoid(-2.25) = 0.09534946
        32'hC00F5C29: sigmoid_out = 32'h3DC50CA7; // -2.24 -> sigmoid(-2.24) = 0.09621554
        32'hC00EB852: sigmoid_out = 32'h3DC6D669; // -2.23 -> sigmoid(-2.23) = 0.09708864
        32'hC00E147B: sigmoid_out = 32'h3DC8A3DE; // -2.22 -> sigmoid(-2.22) = 0.09796880
        32'hC00D70A4: sigmoid_out = 32'h3DCA750E; // -2.21 -> sigmoid(-2.21) = 0.09885607
        32'hC00CCCCD: sigmoid_out = 32'h3DCC49FC; // -2.20 -> sigmoid(-2.20) = 0.09975049
        32'hC00C28F6: sigmoid_out = 32'h3DCE22AF; // -2.19 -> sigmoid(-2.19) = 0.10065209
        32'hC00B851F: sigmoid_out = 32'h3DCFFF2D; // -2.18 -> sigmoid(-2.18) = 0.10156093
        32'hC00AE148: sigmoid_out = 32'h3DD1DF7B; // -2.17 -> sigmoid(-2.17) = 0.10247703
        32'hC00A3D71: sigmoid_out = 32'h3DD3C39E; // -2.16 -> sigmoid(-2.16) = 0.10340045
        32'hC009999A: sigmoid_out = 32'h3DD5AB9C; // -2.15 -> sigmoid(-2.15) = 0.10433122
        32'hC008F5C3: sigmoid_out = 32'h3DD7977A; // -2.14 -> sigmoid(-2.14) = 0.10526939
        32'hC00851EC: sigmoid_out = 32'h3DD9873F; // -2.13 -> sigmoid(-2.13) = 0.10621499
        32'hC007AE14: sigmoid_out = 32'h3DDB7AEF; // -2.12 -> sigmoid(-2.12) = 0.10716807
        32'hC0070A3D: sigmoid_out = 32'h3DDD7290; // -2.11 -> sigmoid(-2.11) = 0.10812867
        32'hC0066666: sigmoid_out = 32'h3DDF6E27; // -2.10 -> sigmoid(-2.10) = 0.10909682
        32'hC005C28F: sigmoid_out = 32'h3DE16DBB; // -2.09 -> sigmoid(-2.09) = 0.11007257
        32'hC0051EB8: sigmoid_out = 32'h3DE37150; // -2.08 -> sigmoid(-2.08) = 0.11105597
        32'hC0047AE1: sigmoid_out = 32'h3DE578EB; // -2.07 -> sigmoid(-2.07) = 0.11204704
        32'hC003D70A: sigmoid_out = 32'h3DE78492; // -2.06 -> sigmoid(-2.06) = 0.11304583
        32'hC0033333: sigmoid_out = 32'h3DE9944B; // -2.05 -> sigmoid(-2.05) = 0.11405238
        32'hC0028F5C: sigmoid_out = 32'h3DEBA81B; // -2.04 -> sigmoid(-2.04) = 0.11506673
        32'hC001EB85: sigmoid_out = 32'h3DEDC007; // -2.03 -> sigmoid(-2.03) = 0.11608892
        32'hC00147AE: sigmoid_out = 32'h3DEFDC15; // -2.02 -> sigmoid(-2.02) = 0.11711899
        32'hC000A3D7: sigmoid_out = 32'h3DF1FC49; // -2.01 -> sigmoid(-2.01) = 0.11815698
        32'hC0000000: sigmoid_out = 32'h3DF420A9; // -2.00 -> sigmoid(-2.00) = 0.11920292
        32'hBFFEB852: sigmoid_out = 32'h3DF6493B; // -1.99 -> sigmoid(-1.99) = 0.12025686
        32'hBFFD70A4: sigmoid_out = 32'h3DF87603; // -1.98 -> sigmoid(-1.98) = 0.12131884
        32'hBFFC28F6: sigmoid_out = 32'h3DFAA706; // -1.97 -> sigmoid(-1.97) = 0.12238889
        32'hBFFAE148: sigmoid_out = 32'h3DFCDC4B; // -1.96 -> sigmoid(-1.96) = 0.12346705
        32'hBFF9999A: sigmoid_out = 32'h3DFF15D5; // -1.95 -> sigmoid(-1.95) = 0.12455336
        32'hBFF851EC: sigmoid_out = 32'h3E00A9D5; // -1.94 -> sigmoid(-1.94) = 0.12564786
        32'hBFF70A3D: sigmoid_out = 32'h3E01CAE7; // -1.93 -> sigmoid(-1.93) = 0.12675058
        32'hBFF5C28F: sigmoid_out = 32'h3E02EE24; // -1.92 -> sigmoid(-1.92) = 0.12786157
        32'hBFF47AE1: sigmoid_out = 32'h3E04138E; // -1.91 -> sigmoid(-1.91) = 0.12898085
        32'hBFF33333: sigmoid_out = 32'h3E053B28; // -1.90 -> sigmoid(-1.90) = 0.13010847
        32'hBFF1EB85: sigmoid_out = 32'h3E0664F3; // -1.89 -> sigmoid(-1.89) = 0.13124447
        32'hBFF0A3D7: sigmoid_out = 32'h3E0790F3; // -1.88 -> sigmoid(-1.88) = 0.13238887
        32'hBFEF5C29: sigmoid_out = 32'h3E08BF29; // -1.87 -> sigmoid(-1.87) = 0.13354172
        32'hBFEE147B: sigmoid_out = 32'h3E09EF99; // -1.86 -> sigmoid(-1.86) = 0.13470305
        32'hBFECCCCD: sigmoid_out = 32'h3E0B2244; // -1.85 -> sigmoid(-1.85) = 0.13587290
        32'hBFEB851F: sigmoid_out = 32'h3E0C572D; // -1.84 -> sigmoid(-1.84) = 0.13705129
        32'hBFEA3D71: sigmoid_out = 32'h3E0D8E55; // -1.83 -> sigmoid(-1.83) = 0.13823827
        32'hBFE8F5C3: sigmoid_out = 32'h3E0EC7C1; // -1.82 -> sigmoid(-1.82) = 0.13943387
        32'hBFE7AE14: sigmoid_out = 32'h3E100371; // -1.81 -> sigmoid(-1.81) = 0.14063813
        32'hBFE66666: sigmoid_out = 32'h3E114168; // -1.80 -> sigmoid(-1.80) = 0.14185106
        32'hBFE51EB8: sigmoid_out = 32'h3E1281A8; // -1.79 -> sigmoid(-1.79) = 0.14307272
        32'hBFE3D70A: sigmoid_out = 32'h3E13C433; // -1.78 -> sigmoid(-1.78) = 0.14430313
        32'hBFE28F5C: sigmoid_out = 32'h3E15090C; // -1.77 -> sigmoid(-1.77) = 0.14554233
        32'hBFE147AE: sigmoid_out = 32'h3E165035; // -1.76 -> sigmoid(-1.76) = 0.14679034
        32'hBFE00000: sigmoid_out = 32'h3E1799AF; // -1.75 -> sigmoid(-1.75) = 0.14804720
        32'hBFDEB852: sigmoid_out = 32'h3E18E57D; // -1.74 -> sigmoid(-1.74) = 0.14931293
        32'hBFDD70A4: sigmoid_out = 32'h3E1A33A1; // -1.73 -> sigmoid(-1.73) = 0.15058758
        32'hBFDC28F6: sigmoid_out = 32'h3E1B841D; // -1.72 -> sigmoid(-1.72) = 0.15187116
        32'hBFDAE148: sigmoid_out = 32'h3E1CD6F3; // -1.71 -> sigmoid(-1.71) = 0.15316372
        32'hBFD9999A: sigmoid_out = 32'h3E1E2C24; // -1.70 -> sigmoid(-1.70) = 0.15446527
        32'hBFD851EC: sigmoid_out = 32'h3E1F83B4; // -1.69 -> sigmoid(-1.69) = 0.15577584
        32'hBFD70A3D: sigmoid_out = 32'h3E20DDA2; // -1.68 -> sigmoid(-1.68) = 0.15709547
        32'hBFD5C28F: sigmoid_out = 32'h3E2239F3; // -1.67 -> sigmoid(-1.67) = 0.15842418
        32'hBFD47AE1: sigmoid_out = 32'h3E2398A6; // -1.66 -> sigmoid(-1.66) = 0.15976200
        32'hBFD33333: sigmoid_out = 32'h3E24F9BF; // -1.65 -> sigmoid(-1.65) = 0.16110895
        32'hBFD1EB85: sigmoid_out = 32'h3E265D3E; // -1.64 -> sigmoid(-1.64) = 0.16246506
        32'hBFD0A3D7: sigmoid_out = 32'h3E27C325; // -1.63 -> sigmoid(-1.63) = 0.16383036
        32'hBFCF5C29: sigmoid_out = 32'h3E292B77; // -1.62 -> sigmoid(-1.62) = 0.16520487
        32'hBFCE147B: sigmoid_out = 32'h3E2A9635; // -1.61 -> sigmoid(-1.61) = 0.16658861
        32'hBFCCCCCD: sigmoid_out = 32'h3E2C035F; // -1.60 -> sigmoid(-1.60) = 0.16798161
        32'hBFCB851F: sigmoid_out = 32'h3E2D72F9; // -1.59 -> sigmoid(-1.59) = 0.16938390
        32'hBFCA3D71: sigmoid_out = 32'h3E2EE503; // -1.58 -> sigmoid(-1.58) = 0.17079548
        32'hBFC8F5C3: sigmoid_out = 32'h3E30597E; // -1.57 -> sigmoid(-1.57) = 0.17221639
        32'hBFC7AE14: sigmoid_out = 32'h3E31D06D; // -1.56 -> sigmoid(-1.56) = 0.17364665
        32'hBFC66666: sigmoid_out = 32'h3E3349D1; // -1.55 -> sigmoid(-1.55) = 0.17508627
        32'hBFC51EB8: sigmoid_out = 32'h3E34C5AA; // -1.54 -> sigmoid(-1.54) = 0.17653527
        32'hBFC3D70A: sigmoid_out = 32'h3E3643FA; // -1.53 -> sigmoid(-1.53) = 0.17799369
        32'hBFC28F5C: sigmoid_out = 32'h3E37C4C3; // -1.52 -> sigmoid(-1.52) = 0.17946152
        32'hBFC147AE: sigmoid_out = 32'h3E394805; // -1.51 -> sigmoid(-1.51) = 0.18093879
        32'hBFC00000: sigmoid_out = 32'h3E3ACDC2; // -1.50 -> sigmoid(-1.50) = 0.18242552
        32'hBFBEB852: sigmoid_out = 32'h3E3C55FA; // -1.49 -> sigmoid(-1.49) = 0.18392173
        32'hBFBD70A4: sigmoid_out = 32'h3E3DE0AF; // -1.48 -> sigmoid(-1.48) = 0.18542742
        32'hBFBC28F6: sigmoid_out = 32'h3E3F6DE2; // -1.47 -> sigmoid(-1.47) = 0.18694261
        32'hBFBAE148: sigmoid_out = 32'h3E40FD94; // -1.46 -> sigmoid(-1.46) = 0.18846733
        32'hBFB9999A: sigmoid_out = 32'h3E428FC5; // -1.45 -> sigmoid(-1.45) = 0.19000157
        32'hBFB851EC: sigmoid_out = 32'h3E442477; // -1.44 -> sigmoid(-1.44) = 0.19154535
        32'hBFB70A3D: sigmoid_out = 32'h3E45BBA9; // -1.43 -> sigmoid(-1.43) = 0.19309868
        32'hBFB5C28F: sigmoid_out = 32'h3E47555E; // -1.42 -> sigmoid(-1.42) = 0.19466158
        32'hBFB47AE1: sigmoid_out = 32'h3E48F195; // -1.41 -> sigmoid(-1.41) = 0.19623406
        32'hBFB33333: sigmoid_out = 32'h3E4A904F; // -1.40 -> sigmoid(-1.40) = 0.19781611
        32'hBFB1EB85: sigmoid_out = 32'h3E4C318C; // -1.39 -> sigmoid(-1.39) = 0.19940776
        32'hBFB0A3D7: sigmoid_out = 32'h3E4DD54E; // -1.38 -> sigmoid(-1.38) = 0.20100900
        32'hBFAF5C29: sigmoid_out = 32'h3E4F7B94; // -1.37 -> sigmoid(-1.37) = 0.20261985
        32'hBFAE147B: sigmoid_out = 32'h3E51245F; // -1.36 -> sigmoid(-1.36) = 0.20424030
        32'hBFACCCCD: sigmoid_out = 32'h3E52CFAF; // -1.35 -> sigmoid(-1.35) = 0.20587037
        32'hBFAB851F: sigmoid_out = 32'h3E547D84; // -1.34 -> sigmoid(-1.34) = 0.20751006
        32'hBFAA3D71: sigmoid_out = 32'h3E562DDF; // -1.33 -> sigmoid(-1.33) = 0.20915937
        32'hBFA8F5C3: sigmoid_out = 32'h3E57E0C0; // -1.32 -> sigmoid(-1.32) = 0.21081829
        32'hBFA7AE14: sigmoid_out = 32'h3E599627; // -1.31 -> sigmoid(-1.31) = 0.21248684
        32'hBFA66666: sigmoid_out = 32'h3E5B4E13; // -1.30 -> sigmoid(-1.30) = 0.21416502
        32'hBFA51EB8: sigmoid_out = 32'h3E5D0885; // -1.29 -> sigmoid(-1.29) = 0.21585281
        32'hBFA3D70A: sigmoid_out = 32'h3E5EC57C; // -1.28 -> sigmoid(-1.28) = 0.21755022
        32'hBFA28F5C: sigmoid_out = 32'h3E6084F9; // -1.27 -> sigmoid(-1.27) = 0.21925725
        32'hBFA147AE: sigmoid_out = 32'h3E6246FB; // -1.26 -> sigmoid(-1.26) = 0.22097389
        32'hBFA00000: sigmoid_out = 32'h3E640B81; // -1.25 -> sigmoid(-1.25) = 0.22270014
        32'hBF9EB852: sigmoid_out = 32'h3E65D28C; // -1.24 -> sigmoid(-1.24) = 0.22443599
        32'hBF9D70A4: sigmoid_out = 32'h3E679C1B; // -1.23 -> sigmoid(-1.23) = 0.22618143
        32'hBF9C28F6: sigmoid_out = 32'h3E69682C; // -1.22 -> sigmoid(-1.22) = 0.22793645
        32'hBF9AE148: sigmoid_out = 32'h3E6B36C1; // -1.21 -> sigmoid(-1.21) = 0.22970105
        32'hBF99999A: sigmoid_out = 32'h3E6D07D7; // -1.20 -> sigmoid(-1.20) = 0.23147522
        32'hBF9851EC: sigmoid_out = 32'h3E6EDB6E; // -1.19 -> sigmoid(-1.19) = 0.23325894
        32'hBF970A3D: sigmoid_out = 32'h3E70B186; // -1.18 -> sigmoid(-1.18) = 0.23505220
        32'hBF95C28F: sigmoid_out = 32'h3E728A1D; // -1.17 -> sigmoid(-1.17) = 0.23685498
        32'hBF947AE1: sigmoid_out = 32'h3E746532; // -1.16 -> sigmoid(-1.16) = 0.23866729
        32'hBF933333: sigmoid_out = 32'h3E7642C5; // -1.15 -> sigmoid(-1.15) = 0.24048908
        32'hBF91EB85: sigmoid_out = 32'h3E7822D4; // -1.14 -> sigmoid(-1.14) = 0.24232036
        32'hBF90A3D7: sigmoid_out = 32'h3E7A055E; // -1.13 -> sigmoid(-1.13) = 0.24416110
        32'hBF8F5C29: sigmoid_out = 32'h3E7BEA62; // -1.12 -> sigmoid(-1.12) = 0.24601128
        32'hBF8E147B: sigmoid_out = 32'h3E7DD1DE; // -1.11 -> sigmoid(-1.11) = 0.24787089
        32'hBF8CCCCD: sigmoid_out = 32'h3E7FBBD1; // -1.10 -> sigmoid(-1.10) = 0.24973989
        32'hBF8B851F: sigmoid_out = 32'h3E80D41C; // -1.09 -> sigmoid(-1.09) = 0.25161828
        32'hBF8A3D71: sigmoid_out = 32'h3E81CB8A; // -1.08 -> sigmoid(-1.08) = 0.25350602
        32'hBF88F5C3: sigmoid_out = 32'h3E82C431; // -1.07 -> sigmoid(-1.07) = 0.25540308
        32'hBF87AE14: sigmoid_out = 32'h3E83BE11; // -1.06 -> sigmoid(-1.06) = 0.25730945
        32'hBF866666: sigmoid_out = 32'h3E84B927; // -1.05 -> sigmoid(-1.05) = 0.25922510
        32'hBF851EB8: sigmoid_out = 32'h3E85B574; // -1.04 -> sigmoid(-1.04) = 0.26114999
        32'hBF83D70A: sigmoid_out = 32'h3E86B2F6; // -1.03 -> sigmoid(-1.03) = 0.26308410
        32'hBF828F5C: sigmoid_out = 32'h3E87B1AC; // -1.02 -> sigmoid(-1.02) = 0.26502740
        32'hBF8147AE: sigmoid_out = 32'h3E88B195; // -1.01 -> sigmoid(-1.01) = 0.26697985
        32'hBF800000: sigmoid_out = 32'h3E89B2B1; // -1.00 -> sigmoid(-1.00) = 0.26894142
        32'hBF7D70A4: sigmoid_out = 32'h3E8AB4FD; // -0.99 -> sigmoid(-0.99) = 0.27091208
        32'hBF7AE148: sigmoid_out = 32'h3E8BB879; // -0.98 -> sigmoid(-0.98) = 0.27289178
        32'hBF7851EC: sigmoid_out = 32'h3E8CBD23; // -0.97 -> sigmoid(-0.97) = 0.27488050
        32'hBF75C28F: sigmoid_out = 32'h3E8DC2FB; // -0.96 -> sigmoid(-0.96) = 0.27687819
        32'hBF733333: sigmoid_out = 32'h3E8EC9FE; // -0.95 -> sigmoid(-0.95) = 0.27888482
        32'hBF70A3D7: sigmoid_out = 32'h3E8FD22B; // -0.94 -> sigmoid(-0.94) = 0.28090034
        32'hBF6E147B: sigmoid_out = 32'h3E90DB82; // -0.93 -> sigmoid(-0.93) = 0.28292471
        32'hBF6B851F: sigmoid_out = 32'h3E91E600; // -0.92 -> sigmoid(-0.92) = 0.28495789
        32'hBF68F5C3: sigmoid_out = 32'h3E92F1A5; // -0.91 -> sigmoid(-0.91) = 0.28699984
        32'hBF666666: sigmoid_out = 32'h3E93FE6D; // -0.90 -> sigmoid(-0.90) = 0.28905050
        32'hBF63D70A: sigmoid_out = 32'h3E950C59; // -0.89 -> sigmoid(-0.89) = 0.29110983
        32'hBF6147AE: sigmoid_out = 32'h3E961B66; // -0.88 -> sigmoid(-0.88) = 0.29317778
        32'hBF5EB852: sigmoid_out = 32'h3E972B92; // -0.87 -> sigmoid(-0.87) = 0.29525430
        32'hBF5C28F6: sigmoid_out = 32'h3E983CDD; // -0.86 -> sigmoid(-0.86) = 0.29733935
        32'hBF59999A: sigmoid_out = 32'h3E994F43; // -0.85 -> sigmoid(-0.85) = 0.29943286
        32'hBF570A3D: sigmoid_out = 32'h3E9A62C4; // -0.84 -> sigmoid(-0.84) = 0.30153478
        32'hBF547AE1: sigmoid_out = 32'h3E9B775E; // -0.83 -> sigmoid(-0.83) = 0.30364507
        32'hBF51EB85: sigmoid_out = 32'h3E9C8D0E; // -0.82 -> sigmoid(-0.82) = 0.30576366
        32'hBF4F5C29: sigmoid_out = 32'h3E9DA3D3; // -0.81 -> sigmoid(-0.81) = 0.30789050
        32'hBF4CCCCD: sigmoid_out = 32'h3E9EBBAA; // -0.80 -> sigmoid(-0.80) = 0.31002552
        32'hBF4A3D71: sigmoid_out = 32'h3E9FD492; // -0.79 -> sigmoid(-0.79) = 0.31216867
        32'hBF47AE14: sigmoid_out = 32'h3EA0EE89; // -0.78 -> sigmoid(-0.78) = 0.31431989
        32'hBF451EB8: sigmoid_out = 32'h3EA2098D; // -0.77 -> sigmoid(-0.77) = 0.31647911
        32'hBF428F5C: sigmoid_out = 32'h3EA3259A; // -0.76 -> sigmoid(-0.76) = 0.31864627
        32'hBF400000: sigmoid_out = 32'h3EA442B1; // -0.75 -> sigmoid(-0.75) = 0.32082130
        32'hBF3D70A4: sigmoid_out = 32'h3EA560CD; // -0.74 -> sigmoid(-0.74) = 0.32300414
        32'hBF3AE148: sigmoid_out = 32'h3EA67FEC; // -0.73 -> sigmoid(-0.73) = 0.32519473
        32'hBF3851EC: sigmoid_out = 32'h3EA7A00E; // -0.72 -> sigmoid(-0.72) = 0.32739298
        32'hBF35C28F: sigmoid_out = 32'h3EA8C12E; // -0.71 -> sigmoid(-0.71) = 0.32959884
        32'hBF333333: sigmoid_out = 32'h3EA9E34B; // -0.70 -> sigmoid(-0.70) = 0.33181223
        32'hBF30A3D7: sigmoid_out = 32'h3EAB0662; // -0.69 -> sigmoid(-0.69) = 0.33403307
        32'hBF2E147B: sigmoid_out = 32'h3EAC2A71; // -0.68 -> sigmoid(-0.68) = 0.33626130
        32'hBF2B851F: sigmoid_out = 32'h3EAD4F75; // -0.67 -> sigmoid(-0.67) = 0.33849684
        32'hBF28F5C3: sigmoid_out = 32'h3EAE756C; // -0.66 -> sigmoid(-0.66) = 0.34073961
        32'hBF266666: sigmoid_out = 32'h3EAF9C53; // -0.65 -> sigmoid(-0.65) = 0.34298954
        32'hBF23D70A: sigmoid_out = 32'h3EB0C428; // -0.64 -> sigmoid(-0.64) = 0.34524654
        32'hBF2147AE: sigmoid_out = 32'h3EB1ECE7; // -0.63 -> sigmoid(-0.63) = 0.34751054
        32'hBF1EB852: sigmoid_out = 32'h3EB3168E; // -0.62 -> sigmoid(-0.62) = 0.34978145
        32'hBF1C28F6: sigmoid_out = 32'h3EB4411A; // -0.61 -> sigmoid(-0.61) = 0.35205920
        32'hBF19999A: sigmoid_out = 32'h3EB56C89; // -0.60 -> sigmoid(-0.60) = 0.35434369
        32'hBF170A3D: sigmoid_out = 32'h3EB698D8; // -0.59 -> sigmoid(-0.59) = 0.35663485
        32'hBF147AE1: sigmoid_out = 32'h3EB7C603; // -0.58 -> sigmoid(-0.58) = 0.35893259
        32'hBF11EB85: sigmoid_out = 32'h3EB8F408; // -0.57 -> sigmoid(-0.57) = 0.36123682
        32'hBF0F5C29: sigmoid_out = 32'h3EBA22E5; // -0.56 -> sigmoid(-0.56) = 0.36354746
        32'hBF0CCCCD: sigmoid_out = 32'h3EBB5294; // -0.55 -> sigmoid(-0.55) = 0.36586441
        32'hBF0A3D71: sigmoid_out = 32'h3EBC8315; // -0.54 -> sigmoid(-0.54) = 0.36818758
        32'hBF07AE14: sigmoid_out = 32'h3EBDB464; // -0.53 -> sigmoid(-0.53) = 0.37051689
        32'hBF051EB8: sigmoid_out = 32'h3EBEE67D; // -0.52 -> sigmoid(-0.52) = 0.37285223
        32'hBF028F5C: sigmoid_out = 32'h3EC0195E; // -0.51 -> sigmoid(-0.51) = 0.37519353
        32'hBF000000: sigmoid_out = 32'h3EC14D03; // -0.50 -> sigmoid(-0.50) = 0.37754067
        32'hBEFAE148: sigmoid_out = 32'h3EC28169; // -0.49 -> sigmoid(-0.49) = 0.37989357
        32'hBEF5C28F: sigmoid_out = 32'h3EC3B68D; // -0.48 -> sigmoid(-0.48) = 0.38225213
        32'hBEF0A3D7: sigmoid_out = 32'h3EC4EC6C; // -0.47 -> sigmoid(-0.47) = 0.38461624
        32'hBEEB851F: sigmoid_out = 32'h3EC62302; // -0.46 -> sigmoid(-0.46) = 0.38698582
        32'hBEE66666: sigmoid_out = 32'h3EC75A4B; // -0.45 -> sigmoid(-0.45) = 0.38936077
        32'hBEE147AE: sigmoid_out = 32'h3EC89246; // -0.44 -> sigmoid(-0.44) = 0.39174097
        32'hBEDC28F6: sigmoid_out = 32'h3EC9CAED; // -0.43 -> sigmoid(-0.43) = 0.39412633
        32'hBED70A3D: sigmoid_out = 32'h3ECB043E; // -0.42 -> sigmoid(-0.42) = 0.39651675
        32'hBED1EB85: sigmoid_out = 32'h3ECC3E36; // -0.41 -> sigmoid(-0.41) = 0.39891212
        32'hBECCCCCD: sigmoid_out = 32'h3ECD78D0; // -0.40 -> sigmoid(-0.40) = 0.40131234
        32'hBEC7AE14: sigmoid_out = 32'h3ECEB409; // -0.39 -> sigmoid(-0.39) = 0.40371730
        32'hBEC28F5C: sigmoid_out = 32'h3ECFEFDD; // -0.38 -> sigmoid(-0.38) = 0.40612690
        32'hBEBD70A4: sigmoid_out = 32'h3ED12C4A; // -0.37 -> sigmoid(-0.37) = 0.40854102
        32'hBEB851EC: sigmoid_out = 32'h3ED2694B; // -0.36 -> sigmoid(-0.36) = 0.41095957
        32'hBEB33333: sigmoid_out = 32'h3ED3A6DC; // -0.35 -> sigmoid(-0.35) = 0.41338242
        32'hBEAE147B: sigmoid_out = 32'h3ED4E4FB; // -0.34 -> sigmoid(-0.34) = 0.41580948
        32'hBEA8F5C3: sigmoid_out = 32'h3ED623A3; // -0.33 -> sigmoid(-0.33) = 0.41824062
        32'hBEA3D70A: sigmoid_out = 32'h3ED762D0; // -0.32 -> sigmoid(-0.32) = 0.42067575
        32'hBE9EB852: sigmoid_out = 32'h3ED8A27F; // -0.31 -> sigmoid(-0.31) = 0.42311474
        32'hBE99999A: sigmoid_out = 32'h3ED9E2AC; // -0.30 -> sigmoid(-0.30) = 0.42555748
        32'hBE947AE1: sigmoid_out = 32'h3EDB2353; // -0.29 -> sigmoid(-0.29) = 0.42800387
        32'hBE8F5C29: sigmoid_out = 32'h3EDC6470; // -0.28 -> sigmoid(-0.28) = 0.43045378
        32'hBE8A3D71: sigmoid_out = 32'h3EDDA600; // -0.27 -> sigmoid(-0.27) = 0.43290710
        32'hBE851EB8: sigmoid_out = 32'h3EDEE7FE; // -0.26 -> sigmoid(-0.26) = 0.43536371
        32'hBE800000: sigmoid_out = 32'h3EE02A67; // -0.25 -> sigmoid(-0.25) = 0.43782350
        32'hBE75C28F: sigmoid_out = 32'h3EE16D36; // -0.24 -> sigmoid(-0.24) = 0.44028635
        32'hBE6B851F: sigmoid_out = 32'h3EE2B069; // -0.23 -> sigmoid(-0.23) = 0.44275215
        32'hBE6147AE: sigmoid_out = 32'h3EE3F3FA; // -0.22 -> sigmoid(-0.22) = 0.44522076
        32'hBE570A3D: sigmoid_out = 32'h3EE537E6; // -0.21 -> sigmoid(-0.21) = 0.44769209
        32'hBE4CCCCD: sigmoid_out = 32'h3EE67C29; // -0.20 -> sigmoid(-0.20) = 0.45016600
        32'hBE428F5C: sigmoid_out = 32'h3EE7C0BE; // -0.19 -> sigmoid(-0.19) = 0.45264238
        32'hBE3851EC: sigmoid_out = 32'h3EE905A2; // -0.18 -> sigmoid(-0.18) = 0.45512111
        32'hBE2E147B: sigmoid_out = 32'h3EEA4AD1; // -0.17 -> sigmoid(-0.17) = 0.45760206
        32'hBE23D70A: sigmoid_out = 32'h3EEB9047; // -0.16 -> sigmoid(-0.16) = 0.46008512
        32'hBE19999A: sigmoid_out = 32'h3EECD5FF; // -0.15 -> sigmoid(-0.15) = 0.46257015
        32'hBE0F5C29: sigmoid_out = 32'h3EEE1BF5; // -0.14 -> sigmoid(-0.14) = 0.46505705
        32'hBE051EB8: sigmoid_out = 32'h3EEF6226; // -0.13 -> sigmoid(-0.13) = 0.46754569
        32'hBDF5C28F: sigmoid_out = 32'h3EF0A88D; // -0.12 -> sigmoid(-0.12) = 0.47003595
        32'hBDE147AE: sigmoid_out = 32'h3EF1EF26; // -0.11 -> sigmoid(-0.11) = 0.47252770
        32'hBDCCCCCD: sigmoid_out = 32'h3EF335EE; // -0.10 -> sigmoid(-0.10) = 0.47502081
        32'hBDB851EC: sigmoid_out = 32'h3EF47CDE; // -0.09 -> sigmoid(-0.09) = 0.47751518
        32'hBDA3D70A: sigmoid_out = 32'h3EF5C3F5; // -0.08 -> sigmoid(-0.08) = 0.48001066
        32'hBD8F5C29: sigmoid_out = 32'h3EF70B2D; // -0.07 -> sigmoid(-0.07) = 0.48250714
        32'hBD75C28F: sigmoid_out = 32'h3EF85282; // -0.06 -> sigmoid(-0.06) = 0.48500450
        32'hBD4CCCCD: sigmoid_out = 32'h3EF999F1; // -0.05 -> sigmoid(-0.05) = 0.48750260
        32'hBD23D70A: sigmoid_out = 32'h3EFAE174; // -0.04 -> sigmoid(-0.04) = 0.49000133
        32'hBCF5C28F: sigmoid_out = 32'h3EFC2909; // -0.03 -> sigmoid(-0.03) = 0.49250056
        32'hBCA3D70A: sigmoid_out = 32'h3EFD70A9; // -0.02 -> sigmoid(-0.02) = 0.49500017
        32'hBC23D70A: sigmoid_out = 32'h3EFEB853; // -0.01 -> sigmoid(-0.01) = 0.49750002
        32'hAA100000: sigmoid_out = 32'h3F000000; // -0.00 -> sigmoid(-0.00) = 0.50000000
        32'h3C23D70A: sigmoid_out = 32'h3F00A3D7; // 0.01 -> sigmoid(0.01) = 0.50249998
        32'h3CA3D70A: sigmoid_out = 32'h3F0147AB; // 0.02 -> sigmoid(0.02) = 0.50499983
        32'h3CF5C28F: sigmoid_out = 32'h3F01EB7C; // 0.03 -> sigmoid(0.03) = 0.50749944
        32'h3D23D70A: sigmoid_out = 32'h3F028F46; // 0.04 -> sigmoid(0.04) = 0.50999867
        32'h3D4CCCCD: sigmoid_out = 32'h3F033308; // 0.05 -> sigmoid(0.05) = 0.51249740
        32'h3D75C28F: sigmoid_out = 32'h3F03D6BF; // 0.06 -> sigmoid(0.06) = 0.51499550
        32'h3D8F5C29: sigmoid_out = 32'h3F047A69; // 0.07 -> sigmoid(0.07) = 0.51749286
        32'h3DA3D70A: sigmoid_out = 32'h3F051E05; // 0.08 -> sigmoid(0.08) = 0.51998934
        32'h3DB851EC: sigmoid_out = 32'h3F05C191; // 0.09 -> sigmoid(0.09) = 0.52248482
        32'h3DCCCCCD: sigmoid_out = 32'h3F066509; // 0.10 -> sigmoid(0.10) = 0.52497919
        32'h3DE147AE: sigmoid_out = 32'h3F07086D; // 0.11 -> sigmoid(0.11) = 0.52747230
        32'h3DF5C28F: sigmoid_out = 32'h3F07ABB9; // 0.12 -> sigmoid(0.12) = 0.52996405
        32'h3E051EB8: sigmoid_out = 32'h3F084EED; // 0.13 -> sigmoid(0.13) = 0.53245431
        32'h3E0F5C29: sigmoid_out = 32'h3F08F205; // 0.14 -> sigmoid(0.14) = 0.53494295
        32'h3E19999A: sigmoid_out = 32'h3F099501; // 0.15 -> sigmoid(0.15) = 0.53742985
        32'h3E23D70A: sigmoid_out = 32'h3F0A37DD; // 0.16 -> sigmoid(0.16) = 0.53991488
        32'h3E2E147B: sigmoid_out = 32'h3F0ADA97; // 0.17 -> sigmoid(0.17) = 0.54239794
        32'h3E3851EC: sigmoid_out = 32'h3F0B7D2F; // 0.18 -> sigmoid(0.18) = 0.54487889
        32'h3E428F5C: sigmoid_out = 32'h3F0C1FA1; // 0.19 -> sigmoid(0.19) = 0.54735762
        32'h3E4CCCCD: sigmoid_out = 32'h3F0CC1EC; // 0.20 -> sigmoid(0.20) = 0.54983400
        32'h3E570A3D: sigmoid_out = 32'h3F0D640D; // 0.21 -> sigmoid(0.21) = 0.55230791
        32'h3E6147AE: sigmoid_out = 32'h3F0E0603; // 0.22 -> sigmoid(0.22) = 0.55477924
        32'h3E6B851F: sigmoid_out = 32'h3F0EA7CC; // 0.23 -> sigmoid(0.23) = 0.55724785
        32'h3E75C28F: sigmoid_out = 32'h3F0F4965; // 0.24 -> sigmoid(0.24) = 0.55971365
        32'h3E800000: sigmoid_out = 32'h3F0FEACD; // 0.25 -> sigmoid(0.25) = 0.56217650
        32'h3E851EB8: sigmoid_out = 32'h3F108C01; // 0.26 -> sigmoid(0.26) = 0.56463629
        32'h3E8A3D71: sigmoid_out = 32'h3F112D00; // 0.27 -> sigmoid(0.27) = 0.56709290
        32'h3E8F5C29: sigmoid_out = 32'h3F11CDC8; // 0.28 -> sigmoid(0.28) = 0.56954622
        32'h3E947AE1: sigmoid_out = 32'h3F126E57; // 0.29 -> sigmoid(0.29) = 0.57199613
        32'h3E99999A: sigmoid_out = 32'h3F130EAA; // 0.30 -> sigmoid(0.30) = 0.57444252
        32'h3E9EB852: sigmoid_out = 32'h3F13AEC1; // 0.31 -> sigmoid(0.31) = 0.57688526
        32'h3EA3D70A: sigmoid_out = 32'h3F144E98; // 0.32 -> sigmoid(0.32) = 0.57932425
        32'h3EA8F5C3: sigmoid_out = 32'h3F14EE2F; // 0.33 -> sigmoid(0.33) = 0.58175938
        32'h3EAE147B: sigmoid_out = 32'h3F158D83; // 0.34 -> sigmoid(0.34) = 0.58419052
        32'h3EB33333: sigmoid_out = 32'h3F162C92; // 0.35 -> sigmoid(0.35) = 0.58661758
        32'h3EB851EC: sigmoid_out = 32'h3F16CB5B; // 0.36 -> sigmoid(0.36) = 0.58904043
        32'h3EBD70A4: sigmoid_out = 32'h3F1769DB; // 0.37 -> sigmoid(0.37) = 0.59145898
        32'h3EC28F5C: sigmoid_out = 32'h3F180811; // 0.38 -> sigmoid(0.38) = 0.59387310
        32'h3EC7AE14: sigmoid_out = 32'h3F18A5FC; // 0.39 -> sigmoid(0.39) = 0.59628270
        32'h3ECCCCCD: sigmoid_out = 32'h3F194398; // 0.40 -> sigmoid(0.40) = 0.59868766
        32'h3ED1EB85: sigmoid_out = 32'h3F19E0E5; // 0.41 -> sigmoid(0.41) = 0.60108788
        32'h3ED70A3D: sigmoid_out = 32'h3F1A7DE1; // 0.42 -> sigmoid(0.42) = 0.60348325
        32'h3EDC28F6: sigmoid_out = 32'h3F1B1A89; // 0.43 -> sigmoid(0.43) = 0.60587367
        32'h3EE147AE: sigmoid_out = 32'h3F1BB6DD; // 0.44 -> sigmoid(0.44) = 0.60825903
        32'h3EE66666: sigmoid_out = 32'h3F1C52DA; // 0.45 -> sigmoid(0.45) = 0.61063923
        32'h3EEB851F: sigmoid_out = 32'h3F1CEE7F; // 0.46 -> sigmoid(0.46) = 0.61301418
        32'h3EF0A3D7: sigmoid_out = 32'h3F1D89CA; // 0.47 -> sigmoid(0.47) = 0.61538376
        32'h3EF5C28F: sigmoid_out = 32'h3F1E24BA; // 0.48 -> sigmoid(0.48) = 0.61774787
        32'h3EFAE148: sigmoid_out = 32'h3F1EBF4C; // 0.49 -> sigmoid(0.49) = 0.62010643
        32'h3F000000: sigmoid_out = 32'h3F1F597F; // 0.50 -> sigmoid(0.50) = 0.62245933
        32'h3F028F5C: sigmoid_out = 32'h3F1FF351; // 0.51 -> sigmoid(0.51) = 0.62480647
        32'h3F051EB8: sigmoid_out = 32'h3F208CC2; // 0.52 -> sigmoid(0.52) = 0.62714777
        32'h3F07AE14: sigmoid_out = 32'h3F2125CE; // 0.53 -> sigmoid(0.53) = 0.62948311
        32'h3F0A3D71: sigmoid_out = 32'h3F21BE75; // 0.54 -> sigmoid(0.54) = 0.63181242
        32'h3F0CCCCD: sigmoid_out = 32'h3F2256B6; // 0.55 -> sigmoid(0.55) = 0.63413559
        32'h3F0F5C29: sigmoid_out = 32'h3F22EE8E; // 0.56 -> sigmoid(0.56) = 0.63645254
        32'h3F11EB85: sigmoid_out = 32'h3F2385FC; // 0.57 -> sigmoid(0.57) = 0.63876318
        32'h3F147AE1: sigmoid_out = 32'h3F241CFE; // 0.58 -> sigmoid(0.58) = 0.64106741
        32'h3F170A3D: sigmoid_out = 32'h3F24B394; // 0.59 -> sigmoid(0.59) = 0.64336515
        32'h3F19999A: sigmoid_out = 32'h3F2549BB; // 0.60 -> sigmoid(0.60) = 0.64565631
        32'h3F1C28F6: sigmoid_out = 32'h3F25DF73; // 0.61 -> sigmoid(0.61) = 0.64794080
        32'h3F1EB852: sigmoid_out = 32'h3F2674B9; // 0.62 -> sigmoid(0.62) = 0.65021855
        32'h3F2147AE: sigmoid_out = 32'h3F27098D; // 0.63 -> sigmoid(0.63) = 0.65248946
        32'h3F23D70A: sigmoid_out = 32'h3F279DEC; // 0.64 -> sigmoid(0.64) = 0.65475346
        32'h3F266666: sigmoid_out = 32'h3F2831D6; // 0.65 -> sigmoid(0.65) = 0.65701046
        32'h3F28F5C3: sigmoid_out = 32'h3F28C54A; // 0.66 -> sigmoid(0.66) = 0.65926039
        32'h3F2B851F: sigmoid_out = 32'h3F295845; // 0.67 -> sigmoid(0.67) = 0.66150316
        32'h3F2E147B: sigmoid_out = 32'h3F29EAC7; // 0.68 -> sigmoid(0.68) = 0.66373870
        32'h3F30A3D7: sigmoid_out = 32'h3F2A7CCF; // 0.69 -> sigmoid(0.69) = 0.66596693
        32'h3F333333: sigmoid_out = 32'h3F2B0E5B; // 0.70 -> sigmoid(0.70) = 0.66818777
        32'h3F35C28F: sigmoid_out = 32'h3F2B9F69; // 0.71 -> sigmoid(0.71) = 0.67040116
        32'h3F3851EC: sigmoid_out = 32'h3F2C2FF9; // 0.72 -> sigmoid(0.72) = 0.67260702
        32'h3F3AE148: sigmoid_out = 32'h3F2CC00A; // 0.73 -> sigmoid(0.73) = 0.67480527
        32'h3F3D70A4: sigmoid_out = 32'h3F2D4F9A; // 0.74 -> sigmoid(0.74) = 0.67699586
        32'h3F400000: sigmoid_out = 32'h3F2DDEA8; // 0.75 -> sigmoid(0.75) = 0.67917870
        32'h3F428F5C: sigmoid_out = 32'h3F2E6D33; // 0.76 -> sigmoid(0.76) = 0.68135373
        32'h3F451EB8: sigmoid_out = 32'h3F2EFB3A; // 0.77 -> sigmoid(0.77) = 0.68352089
        32'h3F47AE14: sigmoid_out = 32'h3F2F88BB; // 0.78 -> sigmoid(0.78) = 0.68568011
        32'h3F4A3D71: sigmoid_out = 32'h3F3015B7; // 0.79 -> sigmoid(0.79) = 0.68783133
        32'h3F4CCCCD: sigmoid_out = 32'h3F30A22B; // 0.80 -> sigmoid(0.80) = 0.68997448
        32'h3F4F5C29: sigmoid_out = 32'h3F312E17; // 0.81 -> sigmoid(0.81) = 0.69210950
        32'h3F51EB85: sigmoid_out = 32'h3F31B979; // 0.82 -> sigmoid(0.82) = 0.69423634
        32'h3F547AE1: sigmoid_out = 32'h3F324451; // 0.83 -> sigmoid(0.83) = 0.69635493
        32'h3F570A3D: sigmoid_out = 32'h3F32CE9E; // 0.84 -> sigmoid(0.84) = 0.69846522
        32'h3F59999A: sigmoid_out = 32'h3F33585E; // 0.85 -> sigmoid(0.85) = 0.70056714
        32'h3F5C28F6: sigmoid_out = 32'h3F33E192; // 0.86 -> sigmoid(0.86) = 0.70266065
        32'h3F5EB852: sigmoid_out = 32'h3F346A37; // 0.87 -> sigmoid(0.87) = 0.70474570
        32'h3F6147AE: sigmoid_out = 32'h3F34F24D; // 0.88 -> sigmoid(0.88) = 0.70682222
        32'h3F63D70A: sigmoid_out = 32'h3F3579D4; // 0.89 -> sigmoid(0.89) = 0.70889017
        32'h3F666666: sigmoid_out = 32'h3F3600C9; // 0.90 -> sigmoid(0.90) = 0.71094950
        32'h3F68F5C3: sigmoid_out = 32'h3F36872E; // 0.91 -> sigmoid(0.91) = 0.71300016
        32'h3F6B851F: sigmoid_out = 32'h3F370D00; // 0.92 -> sigmoid(0.92) = 0.71504211
        32'h3F6E147B: sigmoid_out = 32'h3F37923F; // 0.93 -> sigmoid(0.93) = 0.71707529
        32'h3F70A3D7: sigmoid_out = 32'h3F3816EA; // 0.94 -> sigmoid(0.94) = 0.71909966
        32'h3F733333: sigmoid_out = 32'h3F389B01; // 0.95 -> sigmoid(0.95) = 0.72111518
        32'h3F75C28F: sigmoid_out = 32'h3F391E83; // 0.96 -> sigmoid(0.96) = 0.72312181
        32'h3F7851EC: sigmoid_out = 32'h3F39A16E; // 0.97 -> sigmoid(0.97) = 0.72511950
        32'h3F7AE148: sigmoid_out = 32'h3F3A23C4; // 0.98 -> sigmoid(0.98) = 0.72710822
        32'h3F7D70A4: sigmoid_out = 32'h3F3AA582; // 0.99 -> sigmoid(0.99) = 0.72908792
        32'h3F800000: sigmoid_out = 32'h3F3B26A8; // 1.00 -> sigmoid(1.00) = 0.73105858
        32'h3F8147AE: sigmoid_out = 32'h3F3BA735; // 1.01 -> sigmoid(1.01) = 0.73302015
        32'h3F828F5C: sigmoid_out = 32'h3F3C272A; // 1.02 -> sigmoid(1.02) = 0.73497260
        32'h3F83D70A: sigmoid_out = 32'h3F3CA685; // 1.03 -> sigmoid(1.03) = 0.73691590
        32'h3F851EB8: sigmoid_out = 32'h3F3D2546; // 1.04 -> sigmoid(1.04) = 0.73885001
        32'h3F866666: sigmoid_out = 32'h3F3DA36C; // 1.05 -> sigmoid(1.05) = 0.74077490
        32'h3F87AE14: sigmoid_out = 32'h3F3E20F8; // 1.06 -> sigmoid(1.06) = 0.74269055
        32'h3F88F5C3: sigmoid_out = 32'h3F3E9DE7; // 1.07 -> sigmoid(1.07) = 0.74459692
        32'h3F8A3D71: sigmoid_out = 32'h3F3F1A3B; // 1.08 -> sigmoid(1.08) = 0.74649398
        32'h3F8B851F: sigmoid_out = 32'h3F3F95F2; // 1.09 -> sigmoid(1.09) = 0.74838172
        32'h3F8CCCCD: sigmoid_out = 32'h3F40110C; // 1.10 -> sigmoid(1.10) = 0.75026011
        32'h3F8E147B: sigmoid_out = 32'h3F408B89; // 1.11 -> sigmoid(1.11) = 0.75212911
        32'h3F8F5C29: sigmoid_out = 32'h3F410568; // 1.12 -> sigmoid(1.12) = 0.75398872
        32'h3F90A3D7: sigmoid_out = 32'h3F417EA8; // 1.13 -> sigmoid(1.13) = 0.75583890
        32'h3F91EB85: sigmoid_out = 32'h3F41F74B; // 1.14 -> sigmoid(1.14) = 0.75767964
        32'h3F933333: sigmoid_out = 32'h3F426F4F; // 1.15 -> sigmoid(1.15) = 0.75951092
        32'h3F947AE1: sigmoid_out = 32'h3F42E6B3; // 1.16 -> sigmoid(1.16) = 0.76133271
        32'h3F95C28F: sigmoid_out = 32'h3F435D79; // 1.17 -> sigmoid(1.17) = 0.76314502
        32'h3F970A3D: sigmoid_out = 32'h3F43D39F; // 1.18 -> sigmoid(1.18) = 0.76494780
        32'h3F9851EC: sigmoid_out = 32'h3F444924; // 1.19 -> sigmoid(1.19) = 0.76674106
        32'h3F99999A: sigmoid_out = 32'h3F44BE0A; // 1.20 -> sigmoid(1.20) = 0.76852478
        32'h3F9AE148: sigmoid_out = 32'h3F453250; // 1.21 -> sigmoid(1.21) = 0.77029895
        32'h3F9C28F6: sigmoid_out = 32'h3F45A5F5; // 1.22 -> sigmoid(1.22) = 0.77206355
        32'h3F9D70A4: sigmoid_out = 32'h3F4618F9; // 1.23 -> sigmoid(1.23) = 0.77381857
        32'h3F9EB852: sigmoid_out = 32'h3F468B5D; // 1.24 -> sigmoid(1.24) = 0.77556401
        32'h3FA00000: sigmoid_out = 32'h3F46FD20; // 1.25 -> sigmoid(1.25) = 0.77729986
        32'h3FA147AE: sigmoid_out = 32'h3F476E41; // 1.26 -> sigmoid(1.26) = 0.77902611
        32'h3FA28F5C: sigmoid_out = 32'h3F47DEC2; // 1.27 -> sigmoid(1.27) = 0.78074275
        32'h3FA3D70A: sigmoid_out = 32'h3F484EA1; // 1.28 -> sigmoid(1.28) = 0.78244978
        32'h3FA51EB8: sigmoid_out = 32'h3F48BDDF; // 1.29 -> sigmoid(1.29) = 0.78414719
        32'h3FA66666: sigmoid_out = 32'h3F492C7B; // 1.30 -> sigmoid(1.30) = 0.78583498
        32'h3FA7AE14: sigmoid_out = 32'h3F499A76; // 1.31 -> sigmoid(1.31) = 0.78751316
        32'h3FA8F5C3: sigmoid_out = 32'h3F4A07D0; // 1.32 -> sigmoid(1.32) = 0.78918171
        32'h3FAA3D71: sigmoid_out = 32'h3F4A7488; // 1.33 -> sigmoid(1.33) = 0.79084063
        32'h3FAB851F: sigmoid_out = 32'h3F4AE09F; // 1.34 -> sigmoid(1.34) = 0.79248994
        32'h3FACCCCD: sigmoid_out = 32'h3F4B4C14; // 1.35 -> sigmoid(1.35) = 0.79412963
        32'h3FAE147B: sigmoid_out = 32'h3F4BB6E8; // 1.36 -> sigmoid(1.36) = 0.79575970
        32'h3FAF5C29: sigmoid_out = 32'h3F4C211B; // 1.37 -> sigmoid(1.37) = 0.79738015
        32'h3FB0A3D7: sigmoid_out = 32'h3F4C8AAD; // 1.38 -> sigmoid(1.38) = 0.79899100
        32'h3FB1EB85: sigmoid_out = 32'h3F4CF39D; // 1.39 -> sigmoid(1.39) = 0.80059224
        32'h3FB33333: sigmoid_out = 32'h3F4D5BEC; // 1.40 -> sigmoid(1.40) = 0.80218389
        32'h3FB47AE1: sigmoid_out = 32'h3F4DC39B; // 1.41 -> sigmoid(1.41) = 0.80376594
        32'h3FB5C28F: sigmoid_out = 32'h3F4E2AA9; // 1.42 -> sigmoid(1.42) = 0.80533842
        32'h3FB70A3D: sigmoid_out = 32'h3F4E9116; // 1.43 -> sigmoid(1.43) = 0.80690132
        32'h3FB851EC: sigmoid_out = 32'h3F4EF6E2; // 1.44 -> sigmoid(1.44) = 0.80845465
        32'h3FB9999A: sigmoid_out = 32'h3F4F5C0F; // 1.45 -> sigmoid(1.45) = 0.80999843
        32'h3FBAE148: sigmoid_out = 32'h3F4FC09B; // 1.46 -> sigmoid(1.46) = 0.81153267
        32'h3FBC28F6: sigmoid_out = 32'h3F502487; // 1.47 -> sigmoid(1.47) = 0.81305739
        32'h3FBD70A4: sigmoid_out = 32'h3F5087D4; // 1.48 -> sigmoid(1.48) = 0.81457258
        32'h3FBEB852: sigmoid_out = 32'h3F50EA81; // 1.49 -> sigmoid(1.49) = 0.81607827
        32'h3FC00000: sigmoid_out = 32'h3F514C90; // 1.50 -> sigmoid(1.50) = 0.81757448
        32'h3FC147AE: sigmoid_out = 32'h3F51ADFF; // 1.51 -> sigmoid(1.51) = 0.81906121
        32'h3FC28F5C: sigmoid_out = 32'h3F520ECF; // 1.52 -> sigmoid(1.52) = 0.82053848
        32'h3FC3D70A: sigmoid_out = 32'h3F526F01; // 1.53 -> sigmoid(1.53) = 0.82200631
        32'h3FC51EB8: sigmoid_out = 32'h3F52CE96; // 1.54 -> sigmoid(1.54) = 0.82346473
        32'h3FC66666: sigmoid_out = 32'h3F532D8C; // 1.55 -> sigmoid(1.55) = 0.82491373
        32'h3FC7AE14: sigmoid_out = 32'h3F538BE5; // 1.56 -> sigmoid(1.56) = 0.82635335
        32'h3FC8F5C3: sigmoid_out = 32'h3F53E9A0; // 1.57 -> sigmoid(1.57) = 0.82778361
        32'h3FCA3D71: sigmoid_out = 32'h3F5446BF; // 1.58 -> sigmoid(1.58) = 0.82920452
        32'h3FCB851F: sigmoid_out = 32'h3F54A342; // 1.59 -> sigmoid(1.59) = 0.83061610
        32'h3FCCCCCD: sigmoid_out = 32'h3F54FF28; // 1.60 -> sigmoid(1.60) = 0.83201839
        32'h3FCE147B: sigmoid_out = 32'h3F555A73; // 1.61 -> sigmoid(1.61) = 0.83341139
        32'h3FCF5C29: sigmoid_out = 32'h3F55B522; // 1.62 -> sigmoid(1.62) = 0.83479513
        32'h3FD0A3D7: sigmoid_out = 32'h3F560F37; // 1.63 -> sigmoid(1.63) = 0.83616964
        32'h3FD1EB85: sigmoid_out = 32'h3F5668B1; // 1.64 -> sigmoid(1.64) = 0.83753494
        32'h3FD33333: sigmoid_out = 32'h3F56C190; // 1.65 -> sigmoid(1.65) = 0.83889105
        32'h3FD47AE1: sigmoid_out = 32'h3F5719D6; // 1.66 -> sigmoid(1.66) = 0.84023800
        32'h3FD5C28F: sigmoid_out = 32'h3F577183; // 1.67 -> sigmoid(1.67) = 0.84157582
        32'h3FD70A3D: sigmoid_out = 32'h3F57C897; // 1.68 -> sigmoid(1.68) = 0.84290453
        32'h3FD851EC: sigmoid_out = 32'h3F581F13; // 1.69 -> sigmoid(1.69) = 0.84422416
        32'h3FD9999A: sigmoid_out = 32'h3F5874F7; // 1.70 -> sigmoid(1.70) = 0.84553473
        32'h3FDAE148: sigmoid_out = 32'h3F58CA43; // 1.71 -> sigmoid(1.71) = 0.84683628
        32'h3FDC28F6: sigmoid_out = 32'h3F591EF9; // 1.72 -> sigmoid(1.72) = 0.84812884
        32'h3FDD70A4: sigmoid_out = 32'h3F597318; // 1.73 -> sigmoid(1.73) = 0.84941242
        32'h3FDEB852: sigmoid_out = 32'h3F59C6A1; // 1.74 -> sigmoid(1.74) = 0.85068707
        32'h3FE00000: sigmoid_out = 32'h3F5A1994; // 1.75 -> sigmoid(1.75) = 0.85195280
        32'h3FE147AE: sigmoid_out = 32'h3F5A6BF3; // 1.76 -> sigmoid(1.76) = 0.85320966
        32'h3FE28F5C: sigmoid_out = 32'h3F5ABDBD; // 1.77 -> sigmoid(1.77) = 0.85445767
        32'h3FE3D70A: sigmoid_out = 32'h3F5B0EF3; // 1.78 -> sigmoid(1.78) = 0.85569687
        32'h3FE51EB8: sigmoid_out = 32'h3F5B5F96; // 1.79 -> sigmoid(1.79) = 0.85692728
        32'h3FE66666: sigmoid_out = 32'h3F5BAFA6; // 1.80 -> sigmoid(1.80) = 0.85814894
        32'h3FE7AE14: sigmoid_out = 32'h3F5BFF24; // 1.81 -> sigmoid(1.81) = 0.85936187
        32'h3FE8F5C3: sigmoid_out = 32'h3F5C4E10; // 1.82 -> sigmoid(1.82) = 0.86056613
        32'h3FEA3D71: sigmoid_out = 32'h3F5C9C6B; // 1.83 -> sigmoid(1.83) = 0.86176173
        32'h3FEB851F: sigmoid_out = 32'h3F5CEA35; // 1.84 -> sigmoid(1.84) = 0.86294871
        32'h3FECCCCD: sigmoid_out = 32'h3F5D376F; // 1.85 -> sigmoid(1.85) = 0.86412710
        32'h3FEE147B: sigmoid_out = 32'h3F5D841A; // 1.86 -> sigmoid(1.86) = 0.86529695
        32'h3FEF5C29: sigmoid_out = 32'h3F5DD036; // 1.87 -> sigmoid(1.87) = 0.86645828
        32'h3FF0A3D7: sigmoid_out = 32'h3F5E1BC3; // 1.88 -> sigmoid(1.88) = 0.86761113
        32'h3FF1EB85: sigmoid_out = 32'h3F5E66C3; // 1.89 -> sigmoid(1.89) = 0.86875553
        32'h3FF33333: sigmoid_out = 32'h3F5EB136; // 1.90 -> sigmoid(1.90) = 0.86989153
        32'h3FF47AE1: sigmoid_out = 32'h3F5EFB1C; // 1.91 -> sigmoid(1.91) = 0.87101915
        32'h3FF5C28F: sigmoid_out = 32'h3F5F4477; // 1.92 -> sigmoid(1.92) = 0.87213843
        32'h3FF70A3D: sigmoid_out = 32'h3F5F8D46; // 1.93 -> sigmoid(1.93) = 0.87324942
        32'h3FF851EC: sigmoid_out = 32'h3F5FD58B; // 1.94 -> sigmoid(1.94) = 0.87435214
        32'h3FF9999A: sigmoid_out = 32'h3F601D45; // 1.95 -> sigmoid(1.95) = 0.87544664
        32'h3FFAE148: sigmoid_out = 32'h3F606477; // 1.96 -> sigmoid(1.96) = 0.87653295
        32'h3FFC28F6: sigmoid_out = 32'h3F60AB1F; // 1.97 -> sigmoid(1.97) = 0.87761111
        32'h3FFD70A4: sigmoid_out = 32'h3F60F140; // 1.98 -> sigmoid(1.98) = 0.87868116
        32'h3FFEB852: sigmoid_out = 32'h3F6136D9; // 1.99 -> sigmoid(1.99) = 0.87974314
        32'h40000000: sigmoid_out = 32'h3F617BEB; // 2.00 -> sigmoid(2.00) = 0.88079708
        32'h4000A3D7: sigmoid_out = 32'h3F61C077; // 2.01 -> sigmoid(2.01) = 0.88184302
        32'h400147AE: sigmoid_out = 32'h3F62047D; // 2.02 -> sigmoid(2.02) = 0.88288101
        32'h4001EB85: sigmoid_out = 32'h3F6247FF; // 2.03 -> sigmoid(2.03) = 0.88391108
        32'h40028F5C: sigmoid_out = 32'h3F628AFD; // 2.04 -> sigmoid(2.04) = 0.88493327
        32'h40033333: sigmoid_out = 32'h3F62CD77; // 2.05 -> sigmoid(2.05) = 0.88594762
        32'h4003D70A: sigmoid_out = 32'h3F630F6E; // 2.06 -> sigmoid(2.06) = 0.88695417
        32'h40047AE1: sigmoid_out = 32'h3F6350E3; // 2.07 -> sigmoid(2.07) = 0.88795296
        32'h40051EB8: sigmoid_out = 32'h3F6391D6; // 2.08 -> sigmoid(2.08) = 0.88894403
        32'h4005C28F: sigmoid_out = 32'h3F63D249; // 2.09 -> sigmoid(2.09) = 0.88992743
        32'h40066666: sigmoid_out = 32'h3F64123B; // 2.10 -> sigmoid(2.10) = 0.89090318
        32'h40070A3D: sigmoid_out = 32'h3F6451AE; // 2.11 -> sigmoid(2.11) = 0.89187133
        32'h4007AE14: sigmoid_out = 32'h3F6490A2; // 2.12 -> sigmoid(2.12) = 0.89283193
        32'h400851EC: sigmoid_out = 32'h3F64CF18; // 2.13 -> sigmoid(2.13) = 0.89378501
        32'h4008F5C3: sigmoid_out = 32'h3F650D11; // 2.14 -> sigmoid(2.14) = 0.89473061
        32'h4009999A: sigmoid_out = 32'h3F654A8D; // 2.15 -> sigmoid(2.15) = 0.89566878
        32'h400A3D71: sigmoid_out = 32'h3F65878C; // 2.16 -> sigmoid(2.16) = 0.89659955
        32'h400AE148: sigmoid_out = 32'h3F65C411; // 2.17 -> sigmoid(2.17) = 0.89752297
        32'h400B851F: sigmoid_out = 32'h3F66001A; // 2.18 -> sigmoid(2.18) = 0.89843907
        32'h400C28F6: sigmoid_out = 32'h3F663BAA; // 2.19 -> sigmoid(2.19) = 0.89934791
        32'h400CCCCD: sigmoid_out = 32'h3F6676C0; // 2.20 -> sigmoid(2.20) = 0.90024951
        32'h400D70A4: sigmoid_out = 32'h3F66B15E; // 2.21 -> sigmoid(2.21) = 0.90114393
        32'h400E147B: sigmoid_out = 32'h3F66EB84; // 2.22 -> sigmoid(2.22) = 0.90203120
        32'h400EB852: sigmoid_out = 32'h3F672533; // 2.23 -> sigmoid(2.23) = 0.90291136
        32'h400F5C29: sigmoid_out = 32'h3F675E6B; // 2.24 -> sigmoid(2.24) = 0.90378446
        32'h40100000: sigmoid_out = 32'h3F67972D; // 2.25 -> sigmoid(2.25) = 0.90465054
        32'h4010A3D7: sigmoid_out = 32'h3F67CF7B; // 2.26 -> sigmoid(2.26) = 0.90550963
        32'h401147AE: sigmoid_out = 32'h3F680753; // 2.27 -> sigmoid(2.27) = 0.90636179
        32'h4011EB85: sigmoid_out = 32'h3F683EB9; // 2.28 -> sigmoid(2.28) = 0.90720705
        32'h40128F5C: sigmoid_out = 32'h3F6875AB; // 2.29 -> sigmoid(2.29) = 0.90804545
        32'h40133333: sigmoid_out = 32'h3F68AC2A; // 2.30 -> sigmoid(2.30) = 0.90887704
        32'h4013D70A: sigmoid_out = 32'h3F68E239; // 2.31 -> sigmoid(2.31) = 0.90970186
        32'h40147AE1: sigmoid_out = 32'h3F6917D6; // 2.32 -> sigmoid(2.32) = 0.91051994
        32'h40151EB8: sigmoid_out = 32'h3F694D03; // 2.33 -> sigmoid(2.33) = 0.91133134
        32'h4015C28F: sigmoid_out = 32'h3F6981C0; // 2.34 -> sigmoid(2.34) = 0.91213609
        32'h40166666: sigmoid_out = 32'h3F69B60F; // 2.35 -> sigmoid(2.35) = 0.91293423
        32'h40170A3D: sigmoid_out = 32'h3F69E9EF; // 2.36 -> sigmoid(2.36) = 0.91372581
        32'h4017AE14: sigmoid_out = 32'h3F6A1D62; // 2.37 -> sigmoid(2.37) = 0.91451086
        32'h401851EC: sigmoid_out = 32'h3F6A5069; // 2.38 -> sigmoid(2.38) = 0.91528943
        32'h4018F5C3: sigmoid_out = 32'h3F6A8303; // 2.39 -> sigmoid(2.39) = 0.91606157
        32'h4019999A: sigmoid_out = 32'h3F6AB532; // 2.40 -> sigmoid(2.40) = 0.91682730
        32'h401A3D71: sigmoid_out = 32'h3F6AE6F6; // 2.41 -> sigmoid(2.41) = 0.91758668
        32'h401AE148: sigmoid_out = 32'h3F6B1850; // 2.42 -> sigmoid(2.42) = 0.91833974
        32'h401B851F: sigmoid_out = 32'h3F6B4941; // 2.43 -> sigmoid(2.43) = 0.91908653
        32'h401C28F6: sigmoid_out = 32'h3F6B79CA; // 2.44 -> sigmoid(2.44) = 0.91982709
        32'h401CCCCD: sigmoid_out = 32'h3F6BA9EA; // 2.45 -> sigmoid(2.45) = 0.92056145
        32'h401D70A4: sigmoid_out = 32'h3F6BD9A4; // 2.46 -> sigmoid(2.46) = 0.92128966
        32'h401E147B: sigmoid_out = 32'h3F6C08F7; // 2.47 -> sigmoid(2.47) = 0.92201176
        32'h401EB852: sigmoid_out = 32'h3F6C37E4; // 2.48 -> sigmoid(2.48) = 0.92272780
        32'h401F5C29: sigmoid_out = 32'h3F6C666B; // 2.49 -> sigmoid(2.49) = 0.92343780
        32'h40200000: sigmoid_out = 32'h3F6C948F; // 2.50 -> sigmoid(2.50) = 0.92414182
        32'h4020A3D7: sigmoid_out = 32'h3F6CC24F; // 2.51 -> sigmoid(2.51) = 0.92483989
        32'h402147AE: sigmoid_out = 32'h3F6CEFAB; // 2.52 -> sigmoid(2.52) = 0.92553205
        32'h4021EB85: sigmoid_out = 32'h3F6D1CA5; // 2.53 -> sigmoid(2.53) = 0.92621835
        32'h40228F5C: sigmoid_out = 32'h3F6D493E; // 2.54 -> sigmoid(2.54) = 0.92689883
        32'h40233333: sigmoid_out = 32'h3F6D7575; // 2.55 -> sigmoid(2.55) = 0.92757351
        32'h4023D70A: sigmoid_out = 32'h3F6DA14C; // 2.56 -> sigmoid(2.56) = 0.92824246
        32'h40247AE1: sigmoid_out = 32'h3F6DCCC4; // 2.57 -> sigmoid(2.57) = 0.92890570
        32'h40251EB8: sigmoid_out = 32'h3F6DF7DC; // 2.58 -> sigmoid(2.58) = 0.92956327
        32'h4025C28F: sigmoid_out = 32'h3F6E2296; // 2.59 -> sigmoid(2.59) = 0.93021522
        32'h40266666: sigmoid_out = 32'h3F6E4CF2; // 2.60 -> sigmoid(2.60) = 0.93086158
        32'h40270A3D: sigmoid_out = 32'h3F6E76F1; // 2.61 -> sigmoid(2.61) = 0.93150240
        32'h4027AE14: sigmoid_out = 32'h3F6EA094; // 2.62 -> sigmoid(2.62) = 0.93213771
        32'h402851EC: sigmoid_out = 32'h3F6EC9DB; // 2.63 -> sigmoid(2.63) = 0.93276755
        32'h4028F5C3: sigmoid_out = 32'h3F6EF2C7; // 2.64 -> sigmoid(2.64) = 0.93339196
        32'h4029999A: sigmoid_out = 32'h3F6F1B58; // 2.65 -> sigmoid(2.65) = 0.93401099
        32'h402A3D71: sigmoid_out = 32'h3F6F4390; // 2.66 -> sigmoid(2.66) = 0.93462467
        32'h402AE148: sigmoid_out = 32'h3F6F6B6F; // 2.67 -> sigmoid(2.67) = 0.93523303
        32'h402B851F: sigmoid_out = 32'h3F6F92F5; // 2.68 -> sigmoid(2.68) = 0.93583612
        32'h402C28F6: sigmoid_out = 32'h3F6FBA23; // 2.69 -> sigmoid(2.69) = 0.93643398
        32'h402CCCCD: sigmoid_out = 32'h3F6FE0FA; // 2.70 -> sigmoid(2.70) = 0.93702664
        32'h402D70A4: sigmoid_out = 32'h3F70077B; // 2.71 -> sigmoid(2.71) = 0.93761415
        32'h402E147B: sigmoid_out = 32'h3F702DA6; // 2.72 -> sigmoid(2.72) = 0.93819653
        32'h402EB852: sigmoid_out = 32'h3F70537B; // 2.73 -> sigmoid(2.73) = 0.93877384
        32'h402F5C29: sigmoid_out = 32'h3F7078FC; // 2.74 -> sigmoid(2.74) = 0.93934610
        32'h40300000: sigmoid_out = 32'h3F709E29; // 2.75 -> sigmoid(2.75) = 0.93991335
        32'h4030A3D7: sigmoid_out = 32'h3F70C303; // 2.76 -> sigmoid(2.76) = 0.94047563
        32'h403147AE: sigmoid_out = 32'h3F70E78A; // 2.77 -> sigmoid(2.77) = 0.94103299
        32'h4031EB85: sigmoid_out = 32'h3F710BBE; // 2.78 -> sigmoid(2.78) = 0.94158544
        32'h40328F5C: sigmoid_out = 32'h3F712FA2; // 2.79 -> sigmoid(2.79) = 0.94213304
        32'h40333333: sigmoid_out = 32'h3F715334; // 2.80 -> sigmoid(2.80) = 0.94267582
        32'h4033D70A: sigmoid_out = 32'h3F717676; // 2.81 -> sigmoid(2.81) = 0.94321382
        32'h40347AE1: sigmoid_out = 32'h3F719968; // 2.82 -> sigmoid(2.82) = 0.94374707
        32'h40351EB8: sigmoid_out = 32'h3F71BC0C; // 2.83 -> sigmoid(2.83) = 0.94427560
        32'h4035C28F: sigmoid_out = 32'h3F71DE61; // 2.84 -> sigmoid(2.84) = 0.94479946
        32'h40366666: sigmoid_out = 32'h3F720068; // 2.85 -> sigmoid(2.85) = 0.94531868
        32'h40370A3D: sigmoid_out = 32'h3F722222; // 2.86 -> sigmoid(2.86) = 0.94583330
        32'h4037AE14: sigmoid_out = 32'h3F72438F; // 2.87 -> sigmoid(2.87) = 0.94634335
        32'h403851EC: sigmoid_out = 32'h3F7264B0; // 2.88 -> sigmoid(2.88) = 0.94684886
        32'h4038F5C3: sigmoid_out = 32'h3F728586; // 2.89 -> sigmoid(2.89) = 0.94734988
        32'h4039999A: sigmoid_out = 32'h3F72A610; // 2.90 -> sigmoid(2.90) = 0.94784644
        32'h403A3D71: sigmoid_out = 32'h3F72C651; // 2.91 -> sigmoid(2.91) = 0.94833856
        32'h403AE148: sigmoid_out = 32'h3F72E648; // 2.92 -> sigmoid(2.92) = 0.94882630
        32'h403B851F: sigmoid_out = 32'h3F7305F5; // 2.93 -> sigmoid(2.93) = 0.94930968
        32'h403C28F6: sigmoid_out = 32'h3F73255B; // 2.94 -> sigmoid(2.94) = 0.94978873
        32'h403CCCCD: sigmoid_out = 32'h3F734478; // 2.95 -> sigmoid(2.95) = 0.95026349
        32'h403D70A4: sigmoid_out = 32'h3F73634E; // 2.96 -> sigmoid(2.96) = 0.95073399
        32'h403E147B: sigmoid_out = 32'h3F7381DD; // 2.97 -> sigmoid(2.97) = 0.95120028
        32'h403EB852: sigmoid_out = 32'h3F73A025; // 2.98 -> sigmoid(2.98) = 0.95166237
        32'h403F5C29: sigmoid_out = 32'h3F73BE28; // 2.99 -> sigmoid(2.99) = 0.95212031
        32'h40400000: sigmoid_out = 32'h3F73DBE6; // 3.00 -> sigmoid(3.00) = 0.95257413
        32'h4040A3D7: sigmoid_out = 32'h3F73F95F; // 3.01 -> sigmoid(3.01) = 0.95302385
        32'h404147AE: sigmoid_out = 32'h3F741694; // 3.02 -> sigmoid(3.02) = 0.95346953
        32'h4041EB85: sigmoid_out = 32'h3F743386; // 3.03 -> sigmoid(3.03) = 0.95391117
        32'h40428F5C: sigmoid_out = 32'h3F745034; // 3.04 -> sigmoid(3.04) = 0.95434883
        32'h40433333: sigmoid_out = 32'h3F746CA1; // 3.05 -> sigmoid(3.05) = 0.95478253
        32'h4043D70A: sigmoid_out = 32'h3F7488CB; // 3.06 -> sigmoid(3.06) = 0.95521230
        32'h40447AE1: sigmoid_out = 32'h3F74A4B4; // 3.07 -> sigmoid(3.07) = 0.95563817
        32'h40451EB8: sigmoid_out = 32'h3F74C05C; // 3.08 -> sigmoid(3.08) = 0.95606018
        32'h4045C28F: sigmoid_out = 32'h3F74DBC4; // 3.09 -> sigmoid(3.09) = 0.95647837
        32'h40466666: sigmoid_out = 32'h3F74F6EC; // 3.10 -> sigmoid(3.10) = 0.95689275
        32'h40470A3D: sigmoid_out = 32'h3F7511D5; // 3.11 -> sigmoid(3.11) = 0.95730336
        32'h4047AE14: sigmoid_out = 32'h3F752C7F; // 3.12 -> sigmoid(3.12) = 0.95771023
        32'h404851EC: sigmoid_out = 32'h3F7546EB; // 3.13 -> sigmoid(3.13) = 0.95811339
        32'h4048F5C3: sigmoid_out = 32'h3F75611A; // 3.14 -> sigmoid(3.14) = 0.95851288
        32'h4049999A: sigmoid_out = 32'h3F757B0B; // 3.15 -> sigmoid(3.15) = 0.95890872
        32'h404A3D71: sigmoid_out = 32'h3F7594BF; // 3.16 -> sigmoid(3.16) = 0.95930095
        32'h404AE148: sigmoid_out = 32'h3F75AE37; // 3.17 -> sigmoid(3.17) = 0.95968958
        32'h404B851F: sigmoid_out = 32'h3F75C774; // 3.18 -> sigmoid(3.18) = 0.96007467
        32'h404C28F6: sigmoid_out = 32'h3F75E075; // 3.19 -> sigmoid(3.19) = 0.96045622
        32'h404CCCCD: sigmoid_out = 32'h3F75F93C; // 3.20 -> sigmoid(3.20) = 0.96083428
        32'h404D70A4: sigmoid_out = 32'h3F7611C9; // 3.21 -> sigmoid(3.21) = 0.96120887
        32'h404E147B: sigmoid_out = 32'h3F762A1C; // 3.22 -> sigmoid(3.22) = 0.96158001
        32'h404EB852: sigmoid_out = 32'h3F764235; // 3.23 -> sigmoid(3.23) = 0.96194775
        32'h404F5C29: sigmoid_out = 32'h3F765A16; // 3.24 -> sigmoid(3.24) = 0.96231211
        32'h40500000: sigmoid_out = 32'h3F7671BF; // 3.25 -> sigmoid(3.25) = 0.96267311
        32'h4050A3D7: sigmoid_out = 32'h3F768930; // 3.26 -> sigmoid(3.26) = 0.96303079
        32'h405147AE: sigmoid_out = 32'h3F76A069; // 3.27 -> sigmoid(3.27) = 0.96338517
        32'h4051EB85: sigmoid_out = 32'h3F76B76C; // 3.28 -> sigmoid(3.28) = 0.96373628
        32'h40528F5C: sigmoid_out = 32'h3F76CE38; // 3.29 -> sigmoid(3.29) = 0.96408415
        32'h40533333: sigmoid_out = 32'h3F76E4CE; // 3.30 -> sigmoid(3.30) = 0.96442881
        32'h4053D70A: sigmoid_out = 32'h3F76FB2F; // 3.31 -> sigmoid(3.31) = 0.96477028
        32'h40547AE1: sigmoid_out = 32'h3F77115B; // 3.32 -> sigmoid(3.32) = 0.96510859
        32'h40551EB8: sigmoid_out = 32'h3F772753; // 3.33 -> sigmoid(3.33) = 0.96544377
        32'h4055C28F: sigmoid_out = 32'h3F773D16; // 3.34 -> sigmoid(3.34) = 0.96577584
        32'h40566666: sigmoid_out = 32'h3F7752A6; // 3.35 -> sigmoid(3.35) = 0.96610484
        32'h40570A3D: sigmoid_out = 32'h3F776802; // 3.36 -> sigmoid(3.36) = 0.96643078
        32'h4057AE14: sigmoid_out = 32'h3F777D2B; // 3.37 -> sigmoid(3.37) = 0.96675369
        32'h405851EC: sigmoid_out = 32'h3F779223; // 3.38 -> sigmoid(3.38) = 0.96707361
        32'h4058F5C3: sigmoid_out = 32'h3F77A6E8; // 3.39 -> sigmoid(3.39) = 0.96739054
        32'h4059999A: sigmoid_out = 32'h3F77BB7C; // 3.40 -> sigmoid(3.40) = 0.96770454
        32'h405A3D71: sigmoid_out = 32'h3F77CFDF; // 3.41 -> sigmoid(3.41) = 0.96801560
        32'h405AE148: sigmoid_out = 32'h3F77E411; // 3.42 -> sigmoid(3.42) = 0.96832377
        32'h405B851F: sigmoid_out = 32'h3F77F813; // 3.43 -> sigmoid(3.43) = 0.96862907
        32'h405C28F6: sigmoid_out = 32'h3F780BE5; // 3.44 -> sigmoid(3.44) = 0.96893152
        32'h405CCCCD: sigmoid_out = 32'h3F781F88; // 3.45 -> sigmoid(3.45) = 0.96923114
        32'h405D70A4: sigmoid_out = 32'h3F7832FC; // 3.46 -> sigmoid(3.46) = 0.96952797
        32'h405E147B: sigmoid_out = 32'h3F784641; // 3.47 -> sigmoid(3.47) = 0.96982202
        32'h405EB852: sigmoid_out = 32'h3F785959; // 3.48 -> sigmoid(3.48) = 0.97011332
        32'h405F5C29: sigmoid_out = 32'h3F786C42; // 3.49 -> sigmoid(3.49) = 0.97040190
        32'h40600000: sigmoid_out = 32'h3F787EFE; // 3.50 -> sigmoid(3.50) = 0.97068777
        32'h4060A3D7: sigmoid_out = 32'h3F78918E; // 3.51 -> sigmoid(3.51) = 0.97097096
        32'h406147AE: sigmoid_out = 32'h3F78A3F0; // 3.52 -> sigmoid(3.52) = 0.97125150
        32'h4061EB85: sigmoid_out = 32'h3F78B627; // 3.53 -> sigmoid(3.53) = 0.97152941
        32'h40628F5C: sigmoid_out = 32'h3F78C832; // 3.54 -> sigmoid(3.54) = 0.97180471
        32'h40633333: sigmoid_out = 32'h3F78DA11; // 3.55 -> sigmoid(3.55) = 0.97207743
        32'h4063D70A: sigmoid_out = 32'h3F78EBC5; // 3.56 -> sigmoid(3.56) = 0.97234758
        32'h40647AE1: sigmoid_out = 32'h3F78FD4F; // 3.57 -> sigmoid(3.57) = 0.97261519
        32'h40651EB8: sigmoid_out = 32'h3F790EAF; // 3.58 -> sigmoid(3.58) = 0.97288028
        32'h4065C28F: sigmoid_out = 32'h3F791FE4; // 3.59 -> sigmoid(3.59) = 0.97314288
        32'h40666666: sigmoid_out = 32'h3F7930F0; // 3.60 -> sigmoid(3.60) = 0.97340301
        32'h40670A3D: sigmoid_out = 32'h3F7941D4; // 3.61 -> sigmoid(3.61) = 0.97366068
        32'h4067AE14: sigmoid_out = 32'h3F79528E; // 3.62 -> sigmoid(3.62) = 0.97391592
        32'h406851EC: sigmoid_out = 32'h3F796320; // 3.63 -> sigmoid(3.63) = 0.97416876
        32'h4068F5C3: sigmoid_out = 32'h3F79738A; // 3.64 -> sigmoid(3.64) = 0.97441921
        32'h4069999A: sigmoid_out = 32'h3F7983CC; // 3.65 -> sigmoid(3.65) = 0.97466730
        32'h406A3D71: sigmoid_out = 32'h3F7993E7; // 3.66 -> sigmoid(3.66) = 0.97491304
        32'h406AE148: sigmoid_out = 32'h3F79A3DA; // 3.67 -> sigmoid(3.67) = 0.97515646
        32'h406B851F: sigmoid_out = 32'h3F79B3A8; // 3.68 -> sigmoid(3.68) = 0.97539757
        32'h406C28F6: sigmoid_out = 32'h3F79C34F; // 3.69 -> sigmoid(3.69) = 0.97563641
        32'h406CCCCD: sigmoid_out = 32'h3F79D2D0; // 3.70 -> sigmoid(3.70) = 0.97587298
        32'h406D70A4: sigmoid_out = 32'h3F79E22B; // 3.71 -> sigmoid(3.71) = 0.97610731
        32'h406E147B: sigmoid_out = 32'h3F79F161; // 3.72 -> sigmoid(3.72) = 0.97633942
        32'h406EB852: sigmoid_out = 32'h3F7A0073; // 3.73 -> sigmoid(3.73) = 0.97656933
        32'h406F5C29: sigmoid_out = 32'h3F7A0F5F; // 3.74 -> sigmoid(3.74) = 0.97679706
        32'h40700000: sigmoid_out = 32'h3F7A1E28; // 3.75 -> sigmoid(3.75) = 0.97702263
        32'h4070A3D7: sigmoid_out = 32'h3F7A2CCC; // 3.76 -> sigmoid(3.76) = 0.97724606
        32'h407147AE: sigmoid_out = 32'h3F7A3B4D; // 3.77 -> sigmoid(3.77) = 0.97746736
        32'h4071EB85: sigmoid_out = 32'h3F7A49AB; // 3.78 -> sigmoid(3.78) = 0.97768656
        32'h40728F5C: sigmoid_out = 32'h3F7A57E5; // 3.79 -> sigmoid(3.79) = 0.97790368
        32'h40733333: sigmoid_out = 32'h3F7A65FD; // 3.80 -> sigmoid(3.80) = 0.97811873
        32'h4073D70A: sigmoid_out = 32'h3F7A73F3; // 3.81 -> sigmoid(3.81) = 0.97833173
        32'h40747AE1: sigmoid_out = 32'h3F7A81C6; // 3.82 -> sigmoid(3.82) = 0.97854271
        32'h40751EB8: sigmoid_out = 32'h3F7A8F78; // 3.83 -> sigmoid(3.83) = 0.97875168
        32'h4075C28F: sigmoid_out = 32'h3F7A9D09; // 3.84 -> sigmoid(3.84) = 0.97895865
        32'h40766666: sigmoid_out = 32'h3F7AAA78; // 3.85 -> sigmoid(3.85) = 0.97916366
        32'h40770A3D: sigmoid_out = 32'h3F7AB7C7; // 3.86 -> sigmoid(3.86) = 0.97936670
        32'h4077AE14: sigmoid_out = 32'h3F7AC4F5; // 3.87 -> sigmoid(3.87) = 0.97956781
        32'h407851EC: sigmoid_out = 32'h3F7AD203; // 3.88 -> sigmoid(3.88) = 0.97976700
        32'h4078F5C3: sigmoid_out = 32'h3F7ADEF1; // 3.89 -> sigmoid(3.89) = 0.97996429
        32'h4079999A: sigmoid_out = 32'h3F7AEBBF; // 3.90 -> sigmoid(3.90) = 0.98015969
        32'h407A3D71: sigmoid_out = 32'h3F7AF86E; // 3.91 -> sigmoid(3.91) = 0.98035323
        32'h407AE148: sigmoid_out = 32'h3F7B04FE; // 3.92 -> sigmoid(3.92) = 0.98054492
        32'h407B851F: sigmoid_out = 32'h3F7B116F; // 3.93 -> sigmoid(3.93) = 0.98073477
        32'h407C28F6: sigmoid_out = 32'h3F7B1DC2; // 3.94 -> sigmoid(3.94) = 0.98092280
        32'h407CCCCD: sigmoid_out = 32'h3F7B29F6; // 3.95 -> sigmoid(3.95) = 0.98110904
        32'h407D70A4: sigmoid_out = 32'h3F7B360D; // 3.96 -> sigmoid(3.96) = 0.98129349
        32'h407E147B: sigmoid_out = 32'h3F7B4206; // 3.97 -> sigmoid(3.97) = 0.98147618
        32'h407EB852: sigmoid_out = 32'h3F7B4DE1; // 3.98 -> sigmoid(3.98) = 0.98165711
        32'h407F5C29: sigmoid_out = 32'h3F7B59A0; // 3.99 -> sigmoid(3.99) = 0.98183631
        32'h40800000: sigmoid_out = 32'h3F7B6541; // 4.00 -> sigmoid(4.00) = 0.98201379
        32'h408051EC: sigmoid_out = 32'h3F7B70C7; // 4.01 -> sigmoid(4.01) = 0.98218957
        32'h4080A3D7: sigmoid_out = 32'h3F7B7C2F; // 4.02 -> sigmoid(4.02) = 0.98236366
        32'h4080F5C3: sigmoid_out = 32'h3F7B877C; // 4.03 -> sigmoid(4.03) = 0.98253608
        32'h408147AE: sigmoid_out = 32'h3F7B92AD; // 4.04 -> sigmoid(4.04) = 0.98270684
        32'h4081999A: sigmoid_out = 32'h3F7B9DC2; // 4.05 -> sigmoid(4.05) = 0.98287597
        32'h4081EB85: sigmoid_out = 32'h3F7BA8BD; // 4.06 -> sigmoid(4.06) = 0.98304346
        32'h40823D71: sigmoid_out = 32'h3F7BB39C; // 4.07 -> sigmoid(4.07) = 0.98320935
        32'h40828F5C: sigmoid_out = 32'h3F7BBE60; // 4.08 -> sigmoid(4.08) = 0.98337364
        32'h4082E148: sigmoid_out = 32'h3F7BC90A; // 4.09 -> sigmoid(4.09) = 0.98353636
        32'h40833333: sigmoid_out = 32'h3F7BD399; // 4.10 -> sigmoid(4.10) = 0.98369750
        32'h4083851F: sigmoid_out = 32'h3F7BDE0F; // 4.11 -> sigmoid(4.11) = 0.98385709
        32'h4083D70A: sigmoid_out = 32'h3F7BE86B; // 4.12 -> sigmoid(4.12) = 0.98401515
        32'h408428F6: sigmoid_out = 32'h3F7BF2AD; // 4.13 -> sigmoid(4.13) = 0.98417169
        32'h40847AE1: sigmoid_out = 32'h3F7BFCD6; // 4.14 -> sigmoid(4.14) = 0.98432671
        32'h4084CCCD: sigmoid_out = 32'h3F7C06E6; // 4.15 -> sigmoid(4.15) = 0.98448024
        32'h40851EB8: sigmoid_out = 32'h3F7C10DD; // 4.16 -> sigmoid(4.16) = 0.98463229
        32'h408570A4: sigmoid_out = 32'h3F7C1ABB; // 4.17 -> sigmoid(4.17) = 0.98478288
        32'h4085C28F: sigmoid_out = 32'h3F7C2481; // 4.18 -> sigmoid(4.18) = 0.98493201
        32'h4086147B: sigmoid_out = 32'h3F7C2E2F; // 4.19 -> sigmoid(4.19) = 0.98507970
        32'h40866666: sigmoid_out = 32'h3F7C37C5; // 4.20 -> sigmoid(4.20) = 0.98522597
        32'h4086B852: sigmoid_out = 32'h3F7C4143; // 4.21 -> sigmoid(4.21) = 0.98537082
        32'h40870A3D: sigmoid_out = 32'h3F7C4AAA; // 4.22 -> sigmoid(4.22) = 0.98551428
        32'h40875C29: sigmoid_out = 32'h3F7C53F9; // 4.23 -> sigmoid(4.23) = 0.98565634
        32'h4087AE14: sigmoid_out = 32'h3F7C5D32; // 4.24 -> sigmoid(4.24) = 0.98579704
        32'h40880000: sigmoid_out = 32'h3F7C6653; // 4.25 -> sigmoid(4.25) = 0.98593637
        32'h408851EC: sigmoid_out = 32'h3F7C6F5F; // 4.26 -> sigmoid(4.26) = 0.98607436
        32'h4088A3D7: sigmoid_out = 32'h3F7C7853; // 4.27 -> sigmoid(4.27) = 0.98621101
        32'h4088F5C3: sigmoid_out = 32'h3F7C8132; // 4.28 -> sigmoid(4.28) = 0.98634634
        32'h408947AE: sigmoid_out = 32'h3F7C89FA; // 4.29 -> sigmoid(4.29) = 0.98648036
        32'h4089999A: sigmoid_out = 32'h3F7C92AD; // 4.30 -> sigmoid(4.30) = 0.98661308
        32'h4089EB85: sigmoid_out = 32'h3F7C9B4A; // 4.31 -> sigmoid(4.31) = 0.98674452
        32'h408A3D71: sigmoid_out = 32'h3F7CA3D2; // 4.32 -> sigmoid(4.32) = 0.98687468
        32'h408A8F5C: sigmoid_out = 32'h3F7CAC44; // 4.33 -> sigmoid(4.33) = 0.98700358
        32'h408AE148: sigmoid_out = 32'h3F7CB4A2; // 4.34 -> sigmoid(4.34) = 0.98713124
        32'h408B3333: sigmoid_out = 32'h3F7CBCEB; // 4.35 -> sigmoid(4.35) = 0.98725765
        32'h408B851F: sigmoid_out = 32'h3F7CC51F; // 4.36 -> sigmoid(4.36) = 0.98738284
        32'h408BD70A: sigmoid_out = 32'h3F7CCD3F; // 4.37 -> sigmoid(4.37) = 0.98750681
        32'h408C28F6: sigmoid_out = 32'h3F7CD54B; // 4.38 -> sigmoid(4.38) = 0.98762959
        32'h408C7AE1: sigmoid_out = 32'h3F7CDD43; // 4.39 -> sigmoid(4.39) = 0.98775117
        32'h408CCCCD: sigmoid_out = 32'h3F7CE527; // 4.40 -> sigmoid(4.40) = 0.98787157
        32'h408D1EB8: sigmoid_out = 32'h3F7CECF7; // 4.41 -> sigmoid(4.41) = 0.98799080
        32'h408D70A4: sigmoid_out = 32'h3F7CF4B4; // 4.42 -> sigmoid(4.42) = 0.98810887
        32'h408DC28F: sigmoid_out = 32'h3F7CFC5E; // 4.43 -> sigmoid(4.43) = 0.98822579
        32'h408E147B: sigmoid_out = 32'h3F7D03F4; // 4.44 -> sigmoid(4.44) = 0.98834158
        32'h408E6666: sigmoid_out = 32'h3F7D0B78; // 4.45 -> sigmoid(4.45) = 0.98845625
        32'h408EB852: sigmoid_out = 32'h3F7D12E9; // 4.46 -> sigmoid(4.46) = 0.98856980
        32'h408F0A3D: sigmoid_out = 32'h3F7D1A48; // 4.47 -> sigmoid(4.47) = 0.98868224
        32'h408F5C29: sigmoid_out = 32'h3F7D2194; // 4.48 -> sigmoid(4.48) = 0.98879359
        32'h408FAE14: sigmoid_out = 32'h3F7D28CE; // 4.49 -> sigmoid(4.49) = 0.98890386
        32'h40900000: sigmoid_out = 32'h3F7D2FF6; // 4.50 -> sigmoid(4.50) = 0.98901306
        32'h409051EC: sigmoid_out = 32'h3F7D370C; // 4.51 -> sigmoid(4.51) = 0.98912119
        32'h4090A3D7: sigmoid_out = 32'h3F7D3E10; // 4.52 -> sigmoid(4.52) = 0.98922827
        32'h4090F5C3: sigmoid_out = 32'h3F7D4503; // 4.53 -> sigmoid(4.53) = 0.98933431
        32'h409147AE: sigmoid_out = 32'h3F7D4BE5; // 4.54 -> sigmoid(4.54) = 0.98943931
        32'h4091999A: sigmoid_out = 32'h3F7D52B6; // 4.55 -> sigmoid(4.55) = 0.98954329
        32'h4091EB85: sigmoid_out = 32'h3F7D5975; // 4.56 -> sigmoid(4.56) = 0.98964626
        32'h40923D71: sigmoid_out = 32'h3F7D6024; // 4.57 -> sigmoid(4.57) = 0.98974823
        32'h40928F5C: sigmoid_out = 32'h3F7D66C2; // 4.58 -> sigmoid(4.58) = 0.98984920
        32'h4092E148: sigmoid_out = 32'h3F7D6D4F; // 4.59 -> sigmoid(4.59) = 0.98994919
        32'h40933333: sigmoid_out = 32'h3F7D73CC; // 4.60 -> sigmoid(4.60) = 0.99004820
        32'h4093851F: sigmoid_out = 32'h3F7D7A39; // 4.61 -> sigmoid(4.61) = 0.99014624
        32'h4093D70A: sigmoid_out = 32'h3F7D8096; // 4.62 -> sigmoid(4.62) = 0.99024333
        32'h409428F6: sigmoid_out = 32'h3F7D86E3; // 4.63 -> sigmoid(4.63) = 0.99033948
        32'h40947AE1: sigmoid_out = 32'h3F7D8D21; // 4.64 -> sigmoid(4.64) = 0.99043468
        32'h4094CCCD: sigmoid_out = 32'h3F7D934E; // 4.65 -> sigmoid(4.65) = 0.99052896
        32'h40951EB8: sigmoid_out = 32'h3F7D996C; // 4.66 -> sigmoid(4.66) = 0.99062231
        32'h409570A4: sigmoid_out = 32'h3F7D9F7B; // 4.67 -> sigmoid(4.67) = 0.99071475
        32'h4095C28F: sigmoid_out = 32'h3F7DA57B; // 4.68 -> sigmoid(4.68) = 0.99080629
        32'h4096147B: sigmoid_out = 32'h3F7DAB6C; // 4.69 -> sigmoid(4.69) = 0.99089694
        32'h40966666: sigmoid_out = 32'h3F7DB14E; // 4.70 -> sigmoid(4.70) = 0.99098670
        32'h4096B852: sigmoid_out = 32'h3F7DB721; // 4.71 -> sigmoid(4.71) = 0.99107558
        32'h40970A3D: sigmoid_out = 32'h3F7DBCE6; // 4.72 -> sigmoid(4.72) = 0.99116360
        32'h40975C29: sigmoid_out = 32'h3F7DC29C; // 4.73 -> sigmoid(4.73) = 0.99125075
        32'h4097AE14: sigmoid_out = 32'h3F7DC844; // 4.74 -> sigmoid(4.74) = 0.99133706
        32'h40980000: sigmoid_out = 32'h3F7DCDDE; // 4.75 -> sigmoid(4.75) = 0.99142251
        32'h409851EC: sigmoid_out = 32'h3F7DD369; // 4.76 -> sigmoid(4.76) = 0.99150714
        32'h4098A3D7: sigmoid_out = 32'h3F7DD8E7; // 4.77 -> sigmoid(4.77) = 0.99159093
        32'h4098F5C3: sigmoid_out = 32'h3F7DDE57; // 4.78 -> sigmoid(4.78) = 0.99167391
        32'h409947AE: sigmoid_out = 32'h3F7DE3BA; // 4.79 -> sigmoid(4.79) = 0.99175607
        32'h4099999A: sigmoid_out = 32'h3F7DE90F; // 4.80 -> sigmoid(4.80) = 0.99183743
        32'h4099EB85: sigmoid_out = 32'h3F7DEE56; // 4.81 -> sigmoid(4.81) = 0.99191799
        32'h409A3D71: sigmoid_out = 32'h3F7DF391; // 4.82 -> sigmoid(4.82) = 0.99199777
        32'h409A8F5C: sigmoid_out = 32'h3F7DF8BE; // 4.83 -> sigmoid(4.83) = 0.99207676
        32'h409AE148: sigmoid_out = 32'h3F7DFDDE; // 4.84 -> sigmoid(4.84) = 0.99215498
        32'h409B3333: sigmoid_out = 32'h3F7E02F2; // 4.85 -> sigmoid(4.85) = 0.99223243
        32'h409B851F: sigmoid_out = 32'h3F7E07F9; // 4.86 -> sigmoid(4.86) = 0.99230912
        32'h409BD70A: sigmoid_out = 32'h3F7E0CF3; // 4.87 -> sigmoid(4.87) = 0.99238507
        32'h409C28F6: sigmoid_out = 32'h3F7E11E0; // 4.88 -> sigmoid(4.88) = 0.99246027
        32'h409C7AE1: sigmoid_out = 32'h3F7E16C2; // 4.89 -> sigmoid(4.89) = 0.99253473
        32'h409CCCCD: sigmoid_out = 32'h3F7E1B97; // 4.90 -> sigmoid(4.90) = 0.99260846
        32'h409D1EB8: sigmoid_out = 32'h3F7E205F; // 4.91 -> sigmoid(4.91) = 0.99268147
        32'h409D70A4: sigmoid_out = 32'h3F7E251C; // 4.92 -> sigmoid(4.92) = 0.99275376
        32'h409DC28F: sigmoid_out = 32'h3F7E29CD; // 4.93 -> sigmoid(4.93) = 0.99282534
        32'h409E147B: sigmoid_out = 32'h3F7E2E72; // 4.94 -> sigmoid(4.94) = 0.99289623
        32'h409E6666: sigmoid_out = 32'h3F7E330C; // 4.95 -> sigmoid(4.95) = 0.99296641
        32'h409EB852: sigmoid_out = 32'h3F7E379A; // 4.96 -> sigmoid(4.96) = 0.99303591
        32'h409F0A3D: sigmoid_out = 32'h3F7E3C1D; // 4.97 -> sigmoid(4.97) = 0.99310473
        32'h409F5C29: sigmoid_out = 32'h3F7E4094; // 4.98 -> sigmoid(4.98) = 0.99317287
        32'h409FAE14: sigmoid_out = 32'h3F7E4500; // 4.99 -> sigmoid(4.99) = 0.99324034
        32'h40A00000: sigmoid_out = 32'h3F7E4961; // 5.00 -> sigmoid(5.00) = 0.99330715
        32'h40A051EC: sigmoid_out = 32'h3F7E4DB6; // 5.01 -> sigmoid(5.01) = 0.99337330
        32'h40A0A3D7: sigmoid_out = 32'h3F7E5201; // 5.02 -> sigmoid(5.02) = 0.99343881
        32'h40A0F5C3: sigmoid_out = 32'h3F7E5642; // 5.03 -> sigmoid(5.03) = 0.99350367
        32'h40A147AE: sigmoid_out = 32'h3F7E5A77; // 5.04 -> sigmoid(5.04) = 0.99356789
        32'h40A1999A: sigmoid_out = 32'h3F7E5EA2; // 5.05 -> sigmoid(5.05) = 0.99363148
        32'h40A1EB85: sigmoid_out = 32'h3F7E62C2; // 5.06 -> sigmoid(5.06) = 0.99369445
        32'h40A23D71: sigmoid_out = 32'h3F7E66D9; // 5.07 -> sigmoid(5.07) = 0.99375680
        32'h40A28F5C: sigmoid_out = 32'h3F7E6AE4; // 5.08 -> sigmoid(5.08) = 0.99381854
        32'h40A2E148: sigmoid_out = 32'h3F7E6EE6; // 5.09 -> sigmoid(5.09) = 0.99387967
        32'h40A33333: sigmoid_out = 32'h3F7E72DD; // 5.10 -> sigmoid(5.10) = 0.99394020
        32'h40A3851F: sigmoid_out = 32'h3F7E76CB; // 5.11 -> sigmoid(5.11) = 0.99400013
        32'h40A3D70A: sigmoid_out = 32'h3F7E7AAF; // 5.12 -> sigmoid(5.12) = 0.99405948
        32'h40A428F6: sigmoid_out = 32'h3F7E7E88; // 5.13 -> sigmoid(5.13) = 0.99411824
        32'h40A47AE1: sigmoid_out = 32'h3F7E8259; // 5.14 -> sigmoid(5.14) = 0.99417642
        32'h40A4CCCD: sigmoid_out = 32'h3F7E861F; // 5.15 -> sigmoid(5.15) = 0.99423403
        32'h40A51EB8: sigmoid_out = 32'h3F7E89DC; // 5.16 -> sigmoid(5.16) = 0.99429108
        32'h40A570A4: sigmoid_out = 32'h3F7E8D90; // 5.17 -> sigmoid(5.17) = 0.99434756
        32'h40A5C28F: sigmoid_out = 32'h3F7E913A; // 5.18 -> sigmoid(5.18) = 0.99440349
        32'h40A6147B: sigmoid_out = 32'h3F7E94DB; // 5.19 -> sigmoid(5.19) = 0.99445887
        32'h40A66666: sigmoid_out = 32'h3F7E9873; // 5.20 -> sigmoid(5.20) = 0.99451370
        32'h40A6B852: sigmoid_out = 32'h3F7E9C02; // 5.21 -> sigmoid(5.21) = 0.99456799
        32'h40A70A3D: sigmoid_out = 32'h3F7E9F88; // 5.22 -> sigmoid(5.22) = 0.99462175
        32'h40A75C29: sigmoid_out = 32'h3F7EA305; // 5.23 -> sigmoid(5.23) = 0.99467498
        32'h40A7AE14: sigmoid_out = 32'h3F7EA679; // 5.24 -> sigmoid(5.24) = 0.99472769
        32'h40A80000: sigmoid_out = 32'h3F7EA9E5; // 5.25 -> sigmoid(5.25) = 0.99477987
        32'h40A851EC: sigmoid_out = 32'h3F7EAD48; // 5.26 -> sigmoid(5.26) = 0.99483155
        32'h40A8A3D7: sigmoid_out = 32'h3F7EB0A2; // 5.27 -> sigmoid(5.27) = 0.99488271
        32'h40A8F5C3: sigmoid_out = 32'h3F7EB3F4; // 5.28 -> sigmoid(5.28) = 0.99493337
        32'h40A947AE: sigmoid_out = 32'h3F7EB73E; // 5.29 -> sigmoid(5.29) = 0.99498353
        32'h40A9999A: sigmoid_out = 32'h3F7EBA7F; // 5.30 -> sigmoid(5.30) = 0.99503320
        32'h40A9EB85: sigmoid_out = 32'h3F7EBDB8; // 5.31 -> sigmoid(5.31) = 0.99508238
        32'h40AA3D71: sigmoid_out = 32'h3F7EC0E9; // 5.32 -> sigmoid(5.32) = 0.99513107
        32'h40AA8F5C: sigmoid_out = 32'h3F7EC412; // 5.33 -> sigmoid(5.33) = 0.99517928
        32'h40AAE148: sigmoid_out = 32'h3F7EC733; // 5.34 -> sigmoid(5.34) = 0.99522702
        32'h40AB3333: sigmoid_out = 32'h3F7ECA4C; // 5.35 -> sigmoid(5.35) = 0.99527429
        32'h40AB851F: sigmoid_out = 32'h3F7ECD5D; // 5.36 -> sigmoid(5.36) = 0.99532109
        32'h40ABD70A: sigmoid_out = 32'h3F7ED066; // 5.37 -> sigmoid(5.37) = 0.99536743
        32'h40AC28F6: sigmoid_out = 32'h3F7ED368; // 5.38 -> sigmoid(5.38) = 0.99541331
        32'h40AC7AE1: sigmoid_out = 32'h3F7ED662; // 5.39 -> sigmoid(5.39) = 0.99545874
        32'h40ACCCCD: sigmoid_out = 32'h3F7ED955; // 5.40 -> sigmoid(5.40) = 0.99550373
        32'h40AD1EB8: sigmoid_out = 32'h3F7EDC40; // 5.41 -> sigmoid(5.41) = 0.99554827
        32'h40AD70A4: sigmoid_out = 32'h3F7EDF24; // 5.42 -> sigmoid(5.42) = 0.99559237
        32'h40ADC28F: sigmoid_out = 32'h3F7EE201; // 5.43 -> sigmoid(5.43) = 0.99563603
        32'h40AE147B: sigmoid_out = 32'h3F7EE4D6; // 5.44 -> sigmoid(5.44) = 0.99567927
        32'h40AE6666: sigmoid_out = 32'h3F7EE7A4; // 5.45 -> sigmoid(5.45) = 0.99572207
        32'h40AEB852: sigmoid_out = 32'h3F7EEA6B; // 5.46 -> sigmoid(5.46) = 0.99576446
        32'h40AF0A3D: sigmoid_out = 32'h3F7EED2C; // 5.47 -> sigmoid(5.47) = 0.99580643
        32'h40AF5C29: sigmoid_out = 32'h3F7EEFE5; // 5.48 -> sigmoid(5.48) = 0.99584798
        32'h40AFAE14: sigmoid_out = 32'h3F7EF297; // 5.49 -> sigmoid(5.49) = 0.99588912
        32'h40B00000: sigmoid_out = 32'h3F7EF542; // 5.50 -> sigmoid(5.50) = 0.99592986
        32'h40B051EC: sigmoid_out = 32'h3F7EF7E7; // 5.51 -> sigmoid(5.51) = 0.99597020
        32'h40B0A3D7: sigmoid_out = 32'h3F7EFA85; // 5.52 -> sigmoid(5.52) = 0.99601013
        32'h40B0F5C3: sigmoid_out = 32'h3F7EFD1D; // 5.53 -> sigmoid(5.53) = 0.99604968
        32'h40B147AE: sigmoid_out = 32'h3F7EFFAD; // 5.54 -> sigmoid(5.54) = 0.99608883
        32'h40B1999A: sigmoid_out = 32'h3F7F0238; // 5.55 -> sigmoid(5.55) = 0.99612760
        32'h40B1EB85: sigmoid_out = 32'h3F7F04BC; // 5.56 -> sigmoid(5.56) = 0.99616598
        32'h40B23D71: sigmoid_out = 32'h3F7F0739; // 5.57 -> sigmoid(5.57) = 0.99620398
        32'h40B28F5C: sigmoid_out = 32'h3F7F09B1; // 5.58 -> sigmoid(5.58) = 0.99624161
        32'h40B2E148: sigmoid_out = 32'h3F7F0C22; // 5.59 -> sigmoid(5.59) = 0.99627887
        32'h40B33333: sigmoid_out = 32'h3F7F0E8D; // 5.60 -> sigmoid(5.60) = 0.99631576
        32'h40B3851F: sigmoid_out = 32'h3F7F10F2; // 5.61 -> sigmoid(5.61) = 0.99635229
        32'h40B3D70A: sigmoid_out = 32'h3F7F1350; // 5.62 -> sigmoid(5.62) = 0.99638845
        32'h40B428F6: sigmoid_out = 32'h3F7F15A9; // 5.63 -> sigmoid(5.63) = 0.99642426
        32'h40B47AE1: sigmoid_out = 32'h3F7F17FC; // 5.64 -> sigmoid(5.64) = 0.99645971
        32'h40B4CCCD: sigmoid_out = 32'h3F7F1A49; // 5.65 -> sigmoid(5.65) = 0.99649481
        32'h40B51EB8: sigmoid_out = 32'h3F7F1C90; // 5.66 -> sigmoid(5.66) = 0.99652957
        32'h40B570A4: sigmoid_out = 32'h3F7F1ED1; // 5.67 -> sigmoid(5.67) = 0.99656398
        32'h40B5C28F: sigmoid_out = 32'h3F7F210D; // 5.68 -> sigmoid(5.68) = 0.99659805
        32'h40B6147B: sigmoid_out = 32'h3F7F2343; // 5.69 -> sigmoid(5.69) = 0.99663179
        32'h40B66666: sigmoid_out = 32'h3F7F2573; // 5.70 -> sigmoid(5.70) = 0.99666519
        32'h40B6B852: sigmoid_out = 32'h3F7F279E; // 5.71 -> sigmoid(5.71) = 0.99669827
        32'h40B70A3D: sigmoid_out = 32'h3F7F29C3; // 5.72 -> sigmoid(5.72) = 0.99673101
        32'h40B75C29: sigmoid_out = 32'h3F7F2BE3; // 5.73 -> sigmoid(5.73) = 0.99676343
        32'h40B7AE14: sigmoid_out = 32'h3F7F2DFE; // 5.74 -> sigmoid(5.74) = 0.99679553
        32'h40B80000: sigmoid_out = 32'h3F7F3013; // 5.75 -> sigmoid(5.75) = 0.99682732
        32'h40B851EC: sigmoid_out = 32'h3F7F3223; // 5.76 -> sigmoid(5.76) = 0.99685879
        32'h40B8A3D7: sigmoid_out = 32'h3F7F342E; // 5.77 -> sigmoid(5.77) = 0.99688995
        32'h40B8F5C3: sigmoid_out = 32'h3F7F3634; // 5.78 -> sigmoid(5.78) = 0.99692080
        32'h40B947AE: sigmoid_out = 32'h3F7F3834; // 5.79 -> sigmoid(5.79) = 0.99695134
        32'h40B9999A: sigmoid_out = 32'h3F7F3A2F; // 5.80 -> sigmoid(5.80) = 0.99698158
        32'h40B9EB85: sigmoid_out = 32'h3F7F3C26; // 5.81 -> sigmoid(5.81) = 0.99701153
        32'h40BA3D71: sigmoid_out = 32'h3F7F3E17; // 5.82 -> sigmoid(5.82) = 0.99704118
        32'h40BA8F5C: sigmoid_out = 32'h3F7F4004; // 5.83 -> sigmoid(5.83) = 0.99707053
        32'h40BAE148: sigmoid_out = 32'h3F7F41EB; // 5.84 -> sigmoid(5.84) = 0.99709959
        32'h40BB3333: sigmoid_out = 32'h3F7F43CE; // 5.85 -> sigmoid(5.85) = 0.99712837
        32'h40BB851F: sigmoid_out = 32'h3F7F45AC; // 5.86 -> sigmoid(5.86) = 0.99715686
        32'h40BBD70A: sigmoid_out = 32'h3F7F4785; // 5.87 -> sigmoid(5.87) = 0.99718507
        32'h40BC28F6: sigmoid_out = 32'h3F7F495A; // 5.88 -> sigmoid(5.88) = 0.99721300
        32'h40BC7AE1: sigmoid_out = 32'h3F7F4B2A; // 5.89 -> sigmoid(5.89) = 0.99724066
        32'h40BCCCCD: sigmoid_out = 32'h3F7F4CF5; // 5.90 -> sigmoid(5.90) = 0.99726804
        32'h40BD1EB8: sigmoid_out = 32'h3F7F4EBC; // 5.91 -> sigmoid(5.91) = 0.99729515
        32'h40BD70A4: sigmoid_out = 32'h3F7F507E; // 5.92 -> sigmoid(5.92) = 0.99732199
        32'h40BDC28F: sigmoid_out = 32'h3F7F523C; // 5.93 -> sigmoid(5.93) = 0.99734857
        32'h40BE147B: sigmoid_out = 32'h3F7F53F6; // 5.94 -> sigmoid(5.94) = 0.99737488
        32'h40BE6666: sigmoid_out = 32'h3F7F55AB; // 5.95 -> sigmoid(5.95) = 0.99740093
        32'h40BEB852: sigmoid_out = 32'h3F7F575C; // 5.96 -> sigmoid(5.96) = 0.99742673
        32'h40BF0A3D: sigmoid_out = 32'h3F7F5908; // 5.97 -> sigmoid(5.97) = 0.99745227
        32'h40BF5C29: sigmoid_out = 32'h3F7F5AB0; // 5.98 -> sigmoid(5.98) = 0.99747755
        32'h40BFAE14: sigmoid_out = 32'h3F7F5C54; // 5.99 -> sigmoid(5.99) = 0.99750259
        32'h40C00000: sigmoid_out = 32'h3F7F5DF4; // 6.00 -> sigmoid(6.00) = 0.99752738
    endcase
end



end

endmodule
